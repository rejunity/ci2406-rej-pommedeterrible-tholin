// This is the unpowered netlist.
module wrapped_as1802 (io_oeb,
    rst_n,
    wb_clk_i,
    custom_settings,
    io_in,
    io_out);
 output io_oeb;
 input rst_n;
 input wb_clk_i;
 input [29:0] custom_settings;
 input [35:0] io_in;
 output [35:0] io_out;

 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire \as1802.D[0] ;
 wire \as1802.D[1] ;
 wire \as1802.D[2] ;
 wire \as1802.D[3] ;
 wire \as1802.D[4] ;
 wire \as1802.D[5] ;
 wire \as1802.D[6] ;
 wire \as1802.D[7] ;
 wire \as1802.EF_l[0] ;
 wire \as1802.EF_l[1] ;
 wire \as1802.EF_l[2] ;
 wire \as1802.EF_l[3] ;
 wire \as1802.MHI[0] ;
 wire \as1802.MHI[1] ;
 wire \as1802.MHI[2] ;
 wire \as1802.MHI[3] ;
 wire \as1802.MHI[4] ;
 wire \as1802.MHI[5] ;
 wire \as1802.MHI[6] ;
 wire \as1802.MHI[7] ;
 wire \as1802.MRD ;
 wire \as1802.P[0] ;
 wire \as1802.P[1] ;
 wire \as1802.P[2] ;
 wire \as1802.P[3] ;
 wire \as1802.T[0] ;
 wire \as1802.T[1] ;
 wire \as1802.T[2] ;
 wire \as1802.T[3] ;
 wire \as1802.T[4] ;
 wire \as1802.T[5] ;
 wire \as1802.T[6] ;
 wire \as1802.T[7] ;
 wire \as1802.X[0] ;
 wire \as1802.X[1] ;
 wire \as1802.X[2] ;
 wire \as1802.X[3] ;
 wire \as1802.addr_buff[0] ;
 wire \as1802.addr_buff[10] ;
 wire \as1802.addr_buff[11] ;
 wire \as1802.addr_buff[12] ;
 wire \as1802.addr_buff[13] ;
 wire \as1802.addr_buff[14] ;
 wire \as1802.addr_buff[15] ;
 wire \as1802.addr_buff[1] ;
 wire \as1802.addr_buff[2] ;
 wire \as1802.addr_buff[3] ;
 wire \as1802.addr_buff[4] ;
 wire \as1802.addr_buff[5] ;
 wire \as1802.addr_buff[6] ;
 wire \as1802.addr_buff[7] ;
 wire \as1802.addr_buff[8] ;
 wire \as1802.addr_buff[9] ;
 wire \as1802.cond_inv ;
 wire \as1802.instr_cycle[0] ;
 wire \as1802.instr_cycle[1] ;
 wire \as1802.instr_cycle[2] ;
 wire \as1802.instr_cycle[3] ;
 wire \as1802.instr_latch[0] ;
 wire \as1802.instr_latch[1] ;
 wire \as1802.instr_latch[2] ;
 wire \as1802.instr_latch[4] ;
 wire \as1802.instr_latch[5] ;
 wire \as1802.instr_latch[6] ;
 wire \as1802.instr_latch[7] ;
 wire \as1802.last_hi_addr[0] ;
 wire \as1802.last_hi_addr[1] ;
 wire \as1802.last_hi_addr[2] ;
 wire \as1802.last_hi_addr[3] ;
 wire \as1802.last_hi_addr[4] ;
 wire \as1802.last_hi_addr[5] ;
 wire \as1802.last_hi_addr[6] ;
 wire \as1802.last_hi_addr[7] ;
 wire \as1802.lda ;
 wire \as1802.mem_cycle[0] ;
 wire \as1802.mem_cycle[1] ;
 wire \as1802.mem_cycle[2] ;
 wire \as1802.mem_write ;
 wire \as1802.regs[0][0] ;
 wire \as1802.regs[0][10] ;
 wire \as1802.regs[0][11] ;
 wire \as1802.regs[0][12] ;
 wire \as1802.regs[0][13] ;
 wire \as1802.regs[0][14] ;
 wire \as1802.regs[0][15] ;
 wire \as1802.regs[0][1] ;
 wire \as1802.regs[0][2] ;
 wire \as1802.regs[0][3] ;
 wire \as1802.regs[0][4] ;
 wire \as1802.regs[0][5] ;
 wire \as1802.regs[0][6] ;
 wire \as1802.regs[0][7] ;
 wire \as1802.regs[0][8] ;
 wire \as1802.regs[0][9] ;
 wire \as1802.regs[10][0] ;
 wire \as1802.regs[10][10] ;
 wire \as1802.regs[10][11] ;
 wire \as1802.regs[10][12] ;
 wire \as1802.regs[10][13] ;
 wire \as1802.regs[10][14] ;
 wire \as1802.regs[10][15] ;
 wire \as1802.regs[10][1] ;
 wire \as1802.regs[10][2] ;
 wire \as1802.regs[10][3] ;
 wire \as1802.regs[10][4] ;
 wire \as1802.regs[10][5] ;
 wire \as1802.regs[10][6] ;
 wire \as1802.regs[10][7] ;
 wire \as1802.regs[10][8] ;
 wire \as1802.regs[10][9] ;
 wire \as1802.regs[11][0] ;
 wire \as1802.regs[11][10] ;
 wire \as1802.regs[11][11] ;
 wire \as1802.regs[11][12] ;
 wire \as1802.regs[11][13] ;
 wire \as1802.regs[11][14] ;
 wire \as1802.regs[11][15] ;
 wire \as1802.regs[11][1] ;
 wire \as1802.regs[11][2] ;
 wire \as1802.regs[11][3] ;
 wire \as1802.regs[11][4] ;
 wire \as1802.regs[11][5] ;
 wire \as1802.regs[11][6] ;
 wire \as1802.regs[11][7] ;
 wire \as1802.regs[11][8] ;
 wire \as1802.regs[11][9] ;
 wire \as1802.regs[12][0] ;
 wire \as1802.regs[12][10] ;
 wire \as1802.regs[12][11] ;
 wire \as1802.regs[12][12] ;
 wire \as1802.regs[12][13] ;
 wire \as1802.regs[12][14] ;
 wire \as1802.regs[12][15] ;
 wire \as1802.regs[12][1] ;
 wire \as1802.regs[12][2] ;
 wire \as1802.regs[12][3] ;
 wire \as1802.regs[12][4] ;
 wire \as1802.regs[12][5] ;
 wire \as1802.regs[12][6] ;
 wire \as1802.regs[12][7] ;
 wire \as1802.regs[12][8] ;
 wire \as1802.regs[12][9] ;
 wire \as1802.regs[13][0] ;
 wire \as1802.regs[13][10] ;
 wire \as1802.regs[13][11] ;
 wire \as1802.regs[13][12] ;
 wire \as1802.regs[13][13] ;
 wire \as1802.regs[13][14] ;
 wire \as1802.regs[13][15] ;
 wire \as1802.regs[13][1] ;
 wire \as1802.regs[13][2] ;
 wire \as1802.regs[13][3] ;
 wire \as1802.regs[13][4] ;
 wire \as1802.regs[13][5] ;
 wire \as1802.regs[13][6] ;
 wire \as1802.regs[13][7] ;
 wire \as1802.regs[13][8] ;
 wire \as1802.regs[13][9] ;
 wire \as1802.regs[14][0] ;
 wire \as1802.regs[14][10] ;
 wire \as1802.regs[14][11] ;
 wire \as1802.regs[14][12] ;
 wire \as1802.regs[14][13] ;
 wire \as1802.regs[14][14] ;
 wire \as1802.regs[14][15] ;
 wire \as1802.regs[14][1] ;
 wire \as1802.regs[14][2] ;
 wire \as1802.regs[14][3] ;
 wire \as1802.regs[14][4] ;
 wire \as1802.regs[14][5] ;
 wire \as1802.regs[14][6] ;
 wire \as1802.regs[14][7] ;
 wire \as1802.regs[14][8] ;
 wire \as1802.regs[14][9] ;
 wire \as1802.regs[15][0] ;
 wire \as1802.regs[15][10] ;
 wire \as1802.regs[15][11] ;
 wire \as1802.regs[15][12] ;
 wire \as1802.regs[15][13] ;
 wire \as1802.regs[15][14] ;
 wire \as1802.regs[15][15] ;
 wire \as1802.regs[15][1] ;
 wire \as1802.regs[15][2] ;
 wire \as1802.regs[15][3] ;
 wire \as1802.regs[15][4] ;
 wire \as1802.regs[15][5] ;
 wire \as1802.regs[15][6] ;
 wire \as1802.regs[15][7] ;
 wire \as1802.regs[15][8] ;
 wire \as1802.regs[15][9] ;
 wire \as1802.regs[1][0] ;
 wire \as1802.regs[1][10] ;
 wire \as1802.regs[1][11] ;
 wire \as1802.regs[1][12] ;
 wire \as1802.regs[1][13] ;
 wire \as1802.regs[1][14] ;
 wire \as1802.regs[1][15] ;
 wire \as1802.regs[1][1] ;
 wire \as1802.regs[1][2] ;
 wire \as1802.regs[1][3] ;
 wire \as1802.regs[1][4] ;
 wire \as1802.regs[1][5] ;
 wire \as1802.regs[1][6] ;
 wire \as1802.regs[1][7] ;
 wire \as1802.regs[1][8] ;
 wire \as1802.regs[1][9] ;
 wire \as1802.regs[2][0] ;
 wire \as1802.regs[2][10] ;
 wire \as1802.regs[2][11] ;
 wire \as1802.regs[2][12] ;
 wire \as1802.regs[2][13] ;
 wire \as1802.regs[2][14] ;
 wire \as1802.regs[2][15] ;
 wire \as1802.regs[2][1] ;
 wire \as1802.regs[2][2] ;
 wire \as1802.regs[2][3] ;
 wire \as1802.regs[2][4] ;
 wire \as1802.regs[2][5] ;
 wire \as1802.regs[2][6] ;
 wire \as1802.regs[2][7] ;
 wire \as1802.regs[2][8] ;
 wire \as1802.regs[2][9] ;
 wire \as1802.regs[3][0] ;
 wire \as1802.regs[3][10] ;
 wire \as1802.regs[3][11] ;
 wire \as1802.regs[3][12] ;
 wire \as1802.regs[3][13] ;
 wire \as1802.regs[3][14] ;
 wire \as1802.regs[3][15] ;
 wire \as1802.regs[3][1] ;
 wire \as1802.regs[3][2] ;
 wire \as1802.regs[3][3] ;
 wire \as1802.regs[3][4] ;
 wire \as1802.regs[3][5] ;
 wire \as1802.regs[3][6] ;
 wire \as1802.regs[3][7] ;
 wire \as1802.regs[3][8] ;
 wire \as1802.regs[3][9] ;
 wire \as1802.regs[4][0] ;
 wire \as1802.regs[4][10] ;
 wire \as1802.regs[4][11] ;
 wire \as1802.regs[4][12] ;
 wire \as1802.regs[4][13] ;
 wire \as1802.regs[4][14] ;
 wire \as1802.regs[4][15] ;
 wire \as1802.regs[4][1] ;
 wire \as1802.regs[4][2] ;
 wire \as1802.regs[4][3] ;
 wire \as1802.regs[4][4] ;
 wire \as1802.regs[4][5] ;
 wire \as1802.regs[4][6] ;
 wire \as1802.regs[4][7] ;
 wire \as1802.regs[4][8] ;
 wire \as1802.regs[4][9] ;
 wire \as1802.regs[5][0] ;
 wire \as1802.regs[5][10] ;
 wire \as1802.regs[5][11] ;
 wire \as1802.regs[5][12] ;
 wire \as1802.regs[5][13] ;
 wire \as1802.regs[5][14] ;
 wire \as1802.regs[5][15] ;
 wire \as1802.regs[5][1] ;
 wire \as1802.regs[5][2] ;
 wire \as1802.regs[5][3] ;
 wire \as1802.regs[5][4] ;
 wire \as1802.regs[5][5] ;
 wire \as1802.regs[5][6] ;
 wire \as1802.regs[5][7] ;
 wire \as1802.regs[5][8] ;
 wire \as1802.regs[5][9] ;
 wire \as1802.regs[6][0] ;
 wire \as1802.regs[6][10] ;
 wire \as1802.regs[6][11] ;
 wire \as1802.regs[6][12] ;
 wire \as1802.regs[6][13] ;
 wire \as1802.regs[6][14] ;
 wire \as1802.regs[6][15] ;
 wire \as1802.regs[6][1] ;
 wire \as1802.regs[6][2] ;
 wire \as1802.regs[6][3] ;
 wire \as1802.regs[6][4] ;
 wire \as1802.regs[6][5] ;
 wire \as1802.regs[6][6] ;
 wire \as1802.regs[6][7] ;
 wire \as1802.regs[6][8] ;
 wire \as1802.regs[6][9] ;
 wire \as1802.regs[7][0] ;
 wire \as1802.regs[7][10] ;
 wire \as1802.regs[7][11] ;
 wire \as1802.regs[7][12] ;
 wire \as1802.regs[7][13] ;
 wire \as1802.regs[7][14] ;
 wire \as1802.regs[7][15] ;
 wire \as1802.regs[7][1] ;
 wire \as1802.regs[7][2] ;
 wire \as1802.regs[7][3] ;
 wire \as1802.regs[7][4] ;
 wire \as1802.regs[7][5] ;
 wire \as1802.regs[7][6] ;
 wire \as1802.regs[7][7] ;
 wire \as1802.regs[7][8] ;
 wire \as1802.regs[7][9] ;
 wire \as1802.regs[8][0] ;
 wire \as1802.regs[8][10] ;
 wire \as1802.regs[8][11] ;
 wire \as1802.regs[8][12] ;
 wire \as1802.regs[8][13] ;
 wire \as1802.regs[8][14] ;
 wire \as1802.regs[8][15] ;
 wire \as1802.regs[8][1] ;
 wire \as1802.regs[8][2] ;
 wire \as1802.regs[8][3] ;
 wire \as1802.regs[8][4] ;
 wire \as1802.regs[8][5] ;
 wire \as1802.regs[8][6] ;
 wire \as1802.regs[8][7] ;
 wire \as1802.regs[8][8] ;
 wire \as1802.regs[8][9] ;
 wire \as1802.regs[9][0] ;
 wire \as1802.regs[9][10] ;
 wire \as1802.regs[9][11] ;
 wire \as1802.regs[9][12] ;
 wire \as1802.regs[9][13] ;
 wire \as1802.regs[9][14] ;
 wire \as1802.regs[9][15] ;
 wire \as1802.regs[9][1] ;
 wire \as1802.regs[9][2] ;
 wire \as1802.regs[9][3] ;
 wire \as1802.regs[9][4] ;
 wire \as1802.regs[9][5] ;
 wire \as1802.regs[9][6] ;
 wire \as1802.regs[9][7] ;
 wire \as1802.regs[9][8] ;
 wire \as1802.regs[9][9] ;
 wire \as1802.will_interrupt ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_2379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__B (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A2 (.DIODE(_3488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__B (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__B (.DIODE(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__C (.DIODE(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__B (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__C (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__B (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__B (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__C (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__D (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__C (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__D (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(_3576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1_N (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__S0 (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A1_N (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1_N (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__S (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A1_N (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A1_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1_N (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__C1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__S (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__B (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__S0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__S1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A1_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__C (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__S (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__S0 (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__S0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__S1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A1 (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A1_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__S0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__S1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A1 (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3920__A1_N (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__S (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__S0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__S1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__B (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A_N (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__B (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A_N (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__D (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A2 (.DIODE(_3503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(\as1802.EF_l[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A2 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B2 (.DIODE(\as1802.EF_l[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__C1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A_N (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__B (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__D (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A3 (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A_N (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A2 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__C (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__C1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__C (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__C1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__C (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A (.DIODE(_3488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A2 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B2 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__B (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__C (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A2 (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A0 (.DIODE(\as1802.P[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A0 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A0 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A0 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A0 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A0 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A0 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A0 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A0 (.DIODE(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A1 (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B1 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A1_N (.DIODE(_3438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A2_N (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A1 (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__D (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__C (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A1 (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__C (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A (.DIODE(_3576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A_N (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__S (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A0 (.DIODE(\as1802.P[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__S (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A0 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__B (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A0 (.DIODE(\as1802.P[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__S (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__B1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__S (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__C1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__C (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__B (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__S0 (.DIODE(_0008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__S1 (.DIODE(_0009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A1_N (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A1 (.DIODE(_0010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__B1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A1_N (.DIODE(_0011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__S0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__S1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__C1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__S (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A_N (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A1 (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__B (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__B (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A2 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__C (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__C (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A_N (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A_N (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A_N (.DIODE(_0866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__S0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__S1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__S (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__S0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__S1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__B1 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A1 (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A0 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A (.DIODE(_3437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__B (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A2 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A0 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A1 (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A0 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A2_N (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B2 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__B1 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A0 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__B (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A1_N (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A2_N (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A0 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B1 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A3 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A0 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__S (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__S (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__A (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__B (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__B (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A0 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__A2 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A1 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B1 (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__C (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A2 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A_N (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A1 (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A2 (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__B (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A2 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S0 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__S1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__B (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__C1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A0 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S0 (.DIODE(_0008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__S1 (.DIODE(_0009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__S (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__S1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A1 (.DIODE(_3470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A2 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__B1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__C (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(_3479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A2 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S0 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__S1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__S1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A_N (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A1 (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A2 (.DIODE(_1241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A0 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__S (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__A1 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__C1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A0 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__B (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__S (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__S (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__S (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__B (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S (.DIODE(_1285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__C (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A0 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A0 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A0 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A0 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A0 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S (.DIODE(_1295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__C (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__C (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__B1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__B1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__B (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A0 (.DIODE(_3437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A2 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__C1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__S (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__C1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A2 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A1_N (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__S (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A0 (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__C1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__C1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A0 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__B1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A1_N (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A2_N (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A1 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__C1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__C1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__B2 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B2 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A0 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__S (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__C1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A1 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A1 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A0 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A0 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__B1 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__B (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__C1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__S (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__S (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5056__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__S (.DIODE(_1517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__S (.DIODE(_1527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__S (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__S (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__S (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__S (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__S (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A0 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A0 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A0 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A0 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__S (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A0 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__S (.DIODE(_1572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__S (.DIODE(_1583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__S (.DIODE(_1582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A0 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A0 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A0 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A0 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__S (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A0 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__S (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__C_N (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A0 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A0 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A0 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A0 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A0 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__S (.DIODE(_1613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__S (.DIODE(_1612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__B (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A0 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A0 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A0 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A0 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A0 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__S (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__S (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__S (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__S (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A1 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__C (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A0 (.DIODE(_1332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A0 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A0 (.DIODE(_1401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(_1443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A0 (.DIODE(_1426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A0 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__S (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A0 (.DIODE(_1498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__S (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A0 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A0 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A0 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A0 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__S (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A0 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__S (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__C_N (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A0 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A0 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A0 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A0 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A0 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__S (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__S (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__C (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A0 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A0 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A0 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A0 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A0 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A0 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__S (.DIODE(_1713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A0 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__S (.DIODE(_1712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A3 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__C (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B1 (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A1 (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A1 (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B1 (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__C1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__C1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__C1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A2 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__C1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__C (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__C (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__C (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A2 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__C (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__C (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__D (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__C (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1_N (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A2_N (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__C (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A1 (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A2 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__B (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B1 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__C (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__C (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A2 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__C (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__D (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_3437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B1 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B2 (.DIODE(_3438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__C (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__D (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__C (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__D (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A1 (.DIODE(_3437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B2 (.DIODE(_3438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__C (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__D (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__C (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A (.DIODE(_3510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__C (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__C_N (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__B (.DIODE(_3576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A1 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__C1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__C (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__C (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B2 (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A2 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__B2 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__C1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__C (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1_N (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A (.DIODE(_3488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__B1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A1_N (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__B1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__B2 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B1 (.DIODE(_3510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B2 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__C1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__C (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__D (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A2 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__B1 (.DIODE(_3510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__B1 (.DIODE(_3488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__C1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B1 (.DIODE(_3510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A1 (.DIODE(_3510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A (.DIODE(_3488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__B1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A (.DIODE(_3510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B2 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__C1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__B1 (.DIODE(_3488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__C1 (.DIODE(_2121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__C (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__B1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__C1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__D1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__C_N (.DIODE(_3576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__D1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B (.DIODE(_3527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A2 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A2 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__C1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__B2 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A2 (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A0 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__C1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__C1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A0 (.DIODE(_2347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__C1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A0 (.DIODE(_2355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A0 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__C1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A0 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A0 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__C1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A0 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__S (.DIODE(_2321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A0 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__B2 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A1 (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A0 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A0 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A0 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A2 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B1 (.DIODE(_2417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B2 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A0 (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__C1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A1 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A0 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__C1 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A0 (.DIODE(_1183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__S (.DIODE(_3443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__C1 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A1 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__B2 (.DIODE(_3527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A0 (.DIODE(_1227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__S (.DIODE(_3443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__C1 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A1 (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B2 (.DIODE(_3527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__C1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__S (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A3 (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__C (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A1 (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__C1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__C (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__C1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6227__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__B (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__B (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__B (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A (.DIODE(_3438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__B1 (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__C1 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__B1 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A1 (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A3 (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__C (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__C1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A4 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A1 (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A2 (.DIODE(_3576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A0 (.DIODE(\as1802.P[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A0 (.DIODE(\as1802.P[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A0 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A0 (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A0 (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A (.DIODE(_3432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__C1 (.DIODE(_3550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B2 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A1 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__B2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__B2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__B2 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(_3444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__C (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__B1 (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__C_N (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B1 (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__C_N (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__B1 (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A1 (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A2 (.DIODE(_3623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__S (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A1 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A2 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B2 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A1 (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__C1 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A (.DIODE(_3476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__C1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__C1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A1 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__C1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A1 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__C1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A (.DIODE(_3477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A1 (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__B1 (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__C1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A (.DIODE(_3475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__C1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A (.DIODE(_3437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A1 (.DIODE(_3478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__A2 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A3 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__B1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A3 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__A (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A1 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__C (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__B1 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A1 (.DIODE(_3438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A2 (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__B2 (.DIODE(_3616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__B1 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A1 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__B2 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__C1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__A1 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__B1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__B2 (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__B1_N (.DIODE(_3217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A0 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__S (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__B2 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__B1 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A1 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__B1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A1_N (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A2_N (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__B2 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A1 (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__B1_N (.DIODE(_3247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__A (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__B1 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__B2 (.DIODE(_2005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__A (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__B2 (.DIODE(_3608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__B1_N (.DIODE(_3278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__B1 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__B1 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__B1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A1 (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__C1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__C1 (.DIODE(_3503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__B1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A1 (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__B2 (.DIODE(_3600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__S (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__A (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A1 (.DIODE(_0500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__B2 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A2 (.DIODE(_3592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__B2 (.DIODE(_3436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A1 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__B2 (.DIODE(_3148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__B1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__B1 (.DIODE(_3514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A3 (.DIODE(_3517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A2 (.DIODE(_2715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__B1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__A1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__B1 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__B2 (.DIODE(_0485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__C (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__B (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__S (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__S (.DIODE(_3378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__A1_N (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__C (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__S (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__S (.DIODE(_3404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__A1 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A1 (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__A1 (.DIODE(_1022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__A1 (.DIODE(_0982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A1 (.DIODE(_1117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__A1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A1 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A1 (.DIODE(_1172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__A1 (.DIODE(_1253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__S (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A1 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__S (.DIODE(_3414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__D1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__A3 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A1 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__A1 (.DIODE(net819));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__A1 (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__CLK (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_3503_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_3473_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_3443_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(\as1802.D[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(\as1802.cond_inv ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(_0011_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(_0010_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(_0009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(_0009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(_0008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(_0008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(_0000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_3464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_2321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_2322_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(_3500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(_3527_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold103_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold106_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold117_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold120_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold144_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold146_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold161_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold174_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold180_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold213_A (.DIODE(\as1802.X[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold315_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold500_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold524_A (.DIODE(\as1802.P[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold558_A (.DIODE(\as1802.P[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold591_A (.DIODE(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold592_A (.DIODE(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold599_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold601_A (.DIODE(\as1802.X[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold610_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold615_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold631_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold636_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold637_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold641_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold644_A (.DIODE(\as1802.D[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold647_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold653_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold658_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold660_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold661_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold663_A (.DIODE(\as1802.D[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold70_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold94_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold97_A (.DIODE(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_split26_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_split27_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_split32_A (.DIODE(net143));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_88 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_6 _3630_ (.A(net174),
    .Y(_3432_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(net120),
    .Y(_3433_));
 sky130_fd_sc_hd__inv_2 _3632_ (.A(net128),
    .Y(_3434_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(net129),
    .Y(_3435_));
 sky130_fd_sc_hd__clkinv_4 _3634_ (.A(net131),
    .Y(_3436_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(net133),
    .Y(_3437_));
 sky130_fd_sc_hd__inv_2 _3636_ (.A(net136),
    .Y(_3438_));
 sky130_fd_sc_hd__inv_2 _3637_ (.A(net57),
    .Y(_3439_));
 sky130_fd_sc_hd__inv_2 _3638_ (.A(net827),
    .Y(_3440_));
 sky130_fd_sc_hd__inv_2 _3639_ (.A(net852),
    .Y(_3441_));
 sky130_fd_sc_hd__inv_6 _3640_ (.A(net163),
    .Y(_3442_));
 sky130_fd_sc_hd__inv_2 _3641_ (.A(net164),
    .Y(_3443_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(net315),
    .Y(_3444_));
 sky130_fd_sc_hd__inv_2 _3643_ (.A(net338),
    .Y(_3445_));
 sky130_fd_sc_hd__inv_2 _3644_ (.A(net377),
    .Y(_3446_));
 sky130_fd_sc_hd__inv_2 _3645_ (.A(net306),
    .Y(_3447_));
 sky130_fd_sc_hd__inv_2 _3646_ (.A(net369),
    .Y(_3448_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(net298),
    .Y(_3449_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(net373),
    .Y(_3450_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(net282),
    .Y(_3451_));
 sky130_fd_sc_hd__inv_2 _3650_ (.A(net461),
    .Y(_3452_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(net302),
    .Y(_3453_));
 sky130_fd_sc_hd__inv_2 _3652_ (.A(net371),
    .Y(_3454_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(net290),
    .Y(_3455_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(net356),
    .Y(_3456_));
 sky130_fd_sc_hd__inv_2 _3655_ (.A(net843),
    .Y(_3457_));
 sky130_fd_sc_hd__inv_2 _3656_ (.A(net375),
    .Y(_3458_));
 sky130_fd_sc_hd__inv_2 _3657_ (.A(\as1802.MHI[4] ),
    .Y(_3459_));
 sky130_fd_sc_hd__inv_2 _3658_ (.A(\as1802.MHI[2] ),
    .Y(_3460_));
 sky130_fd_sc_hd__inv_2 _3659_ (.A(\as1802.MHI[1] ),
    .Y(_3461_));
 sky130_fd_sc_hd__inv_2 _3660_ (.A(\as1802.MHI[0] ),
    .Y(_3462_));
 sky130_fd_sc_hd__inv_2 _3661_ (.A(net171),
    .Y(_3463_));
 sky130_fd_sc_hd__inv_2 _3662_ (.A(net212),
    .Y(_3464_));
 sky130_fd_sc_hd__inv_2 _3663_ (.A(net839),
    .Y(_3465_));
 sky130_fd_sc_hd__inv_2 _3664_ (.A(net185),
    .Y(_3466_));
 sky130_fd_sc_hd__inv_2 _3665_ (.A(_0003_),
    .Y(_3467_));
 sky130_fd_sc_hd__inv_2 _3666_ (.A(net18),
    .Y(_3468_));
 sky130_fd_sc_hd__inv_2 _3667_ (.A(net176),
    .Y(_3469_));
 sky130_fd_sc_hd__inv_8 _3668_ (.A(net175),
    .Y(_3470_));
 sky130_fd_sc_hd__inv_2 _3669_ (.A(net158),
    .Y(_3471_));
 sky130_fd_sc_hd__inv_2 _3670_ (.A(net155),
    .Y(_3472_));
 sky130_fd_sc_hd__inv_2 _3671_ (.A(net153),
    .Y(_3473_));
 sky130_fd_sc_hd__inv_2 _3672_ (.A(net151),
    .Y(_3474_));
 sky130_fd_sc_hd__inv_6 _3673_ (.A(net147),
    .Y(_3475_));
 sky130_fd_sc_hd__inv_4 _3674_ (.A(net244),
    .Y(_3476_));
 sky130_fd_sc_hd__inv_2 _3675_ (.A(net141),
    .Y(_3477_));
 sky130_fd_sc_hd__inv_6 _3676_ (.A(net139),
    .Y(_3478_));
 sky130_fd_sc_hd__inv_2 _3677_ (.A(net7),
    .Y(_3479_));
 sky130_fd_sc_hd__inv_2 _3678_ (.A(net40),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _3679_ (.A(net41),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _3680_ (.A(net42),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _3681_ (.A(net43),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _3682_ (.A(net288),
    .Y(_3480_));
 sky130_fd_sc_hd__nor2_1 _3683_ (.A(net843),
    .B(net352),
    .Y(_3481_));
 sky130_fd_sc_hd__and2_1 _3684_ (.A(_3456_),
    .B(_3481_),
    .X(_3482_));
 sky130_fd_sc_hd__nand2_1 _3685_ (.A(_3456_),
    .B(_3481_),
    .Y(_3483_));
 sky130_fd_sc_hd__nor2_2 _3686_ (.A(_3440_),
    .B(\as1802.instr_latch[6] ),
    .Y(_3484_));
 sky130_fd_sc_hd__or2_4 _3687_ (.A(_3440_),
    .B(\as1802.instr_latch[6] ),
    .X(_3485_));
 sky130_fd_sc_hd__nor2_2 _3688_ (.A(_3441_),
    .B(_3485_),
    .Y(_3486_));
 sky130_fd_sc_hd__nand2_1 _3689_ (.A(net852),
    .B(_3484_),
    .Y(_3487_));
 sky130_fd_sc_hd__nor2_4 _3690_ (.A(net163),
    .B(_3487_),
    .Y(_3488_));
 sky130_fd_sc_hd__nand2_4 _3691_ (.A(_3442_),
    .B(_3486_),
    .Y(_3489_));
 sky130_fd_sc_hd__a21oi_1 _3692_ (.A1(net161),
    .A2(_3488_),
    .B1(net103),
    .Y(_3490_));
 sky130_fd_sc_hd__nor2_1 _3693_ (.A(_3464_),
    .B(_3490_),
    .Y(_3491_));
 sky130_fd_sc_hd__nor2_1 _3694_ (.A(\as1802.instr_latch[5] ),
    .B(net163),
    .Y(_3492_));
 sky130_fd_sc_hd__or2_2 _3695_ (.A(\as1802.instr_latch[5] ),
    .B(net163),
    .X(_3493_));
 sky130_fd_sc_hd__and2_1 _3696_ (.A(\as1802.instr_latch[7] ),
    .B(\as1802.instr_latch[6] ),
    .X(_3494_));
 sky130_fd_sc_hd__nand2_1 _3697_ (.A(\as1802.instr_latch[7] ),
    .B(\as1802.instr_latch[6] ),
    .Y(_3495_));
 sky130_fd_sc_hd__nor2_4 _3698_ (.A(_3493_),
    .B(_3495_),
    .Y(_3496_));
 sky130_fd_sc_hd__or3_4 _3699_ (.A(\as1802.instr_latch[7] ),
    .B(\as1802.instr_latch[6] ),
    .C(_3441_),
    .X(_3497_));
 sky130_fd_sc_hd__nor2_4 _3700_ (.A(net163),
    .B(_3497_),
    .Y(_3498_));
 sky130_fd_sc_hd__or2_1 _3701_ (.A(net163),
    .B(_3497_),
    .X(_3499_));
 sky130_fd_sc_hd__a21oi_4 _3702_ (.A1(net161),
    .A2(_3498_),
    .B1(_3496_),
    .Y(_3500_));
 sky130_fd_sc_hd__a21o_2 _3703_ (.A1(net161),
    .A2(_3498_),
    .B1(_3496_),
    .X(_3501_));
 sky130_fd_sc_hd__nor2_1 _3704_ (.A(net169),
    .B(net810),
    .Y(_3502_));
 sky130_fd_sc_hd__and2_2 _3705_ (.A(net167),
    .B(_3502_),
    .X(_3503_));
 sky130_fd_sc_hd__nand2_2 _3706_ (.A(net167),
    .B(_3502_),
    .Y(_3504_));
 sky130_fd_sc_hd__nand2_1 _3707_ (.A(net119),
    .B(net101),
    .Y(_3505_));
 sky130_fd_sc_hd__nor2_1 _3708_ (.A(net164),
    .B(_3505_),
    .Y(_3506_));
 sky130_fd_sc_hd__or2_1 _3709_ (.A(net95),
    .B(_3506_),
    .X(_3507_));
 sky130_fd_sc_hd__nor2_2 _3710_ (.A(net169),
    .B(_3444_),
    .Y(_3508_));
 sky130_fd_sc_hd__and2_1 _3711_ (.A(net168),
    .B(_3508_),
    .X(_3509_));
 sky130_fd_sc_hd__nand2_2 _3712_ (.A(net168),
    .B(_3508_),
    .Y(_3510_));
 sky130_fd_sc_hd__and2_2 _3713_ (.A(net169),
    .B(\as1802.instr_latch[0] ),
    .X(_3511_));
 sky130_fd_sc_hd__nand2_4 _3714_ (.A(net169),
    .B(net315),
    .Y(_3512_));
 sky130_fd_sc_hd__and3_4 _3715_ (.A(net167),
    .B(net169),
    .C(\as1802.instr_latch[0] ),
    .X(_3513_));
 sky130_fd_sc_hd__nand2_4 _3716_ (.A(net167),
    .B(_3511_),
    .Y(_3514_));
 sky130_fd_sc_hd__and2_1 _3717_ (.A(net169),
    .B(_3444_),
    .X(_3515_));
 sky130_fd_sc_hd__nand2_1 _3718_ (.A(net169),
    .B(_3444_),
    .Y(_3516_));
 sky130_fd_sc_hd__and3_4 _3719_ (.A(net168),
    .B(net170),
    .C(_3444_),
    .X(_3517_));
 sky130_fd_sc_hd__o21ai_2 _3720_ (.A1(net170),
    .A2(net810),
    .B1(net167),
    .Y(_3518_));
 sky130_fd_sc_hd__nand2_1 _3721_ (.A(net164),
    .B(_3502_),
    .Y(_3519_));
 sky130_fd_sc_hd__a21oi_4 _3722_ (.A1(_3518_),
    .A2(_3519_),
    .B1(net161),
    .Y(_3520_));
 sky130_fd_sc_hd__nor2_4 _3723_ (.A(_3507_),
    .B(_3520_),
    .Y(_3521_));
 sky130_fd_sc_hd__or2_1 _3724_ (.A(_3507_),
    .B(_3520_),
    .X(_3522_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(_3440_),
    .B(net809),
    .Y(_3523_));
 sky130_fd_sc_hd__or3_4 _3726_ (.A(\as1802.instr_latch[5] ),
    .B(_3442_),
    .C(_3523_),
    .X(_3524_));
 sky130_fd_sc_hd__or3_4 _3727_ (.A(_3441_),
    .B(net163),
    .C(_3523_),
    .X(_3525_));
 sky130_fd_sc_hd__and2_4 _3728_ (.A(_3524_),
    .B(_3525_),
    .X(_3526_));
 sky130_fd_sc_hd__nor2_4 _3729_ (.A(_3442_),
    .B(_3497_),
    .Y(_3527_));
 sky130_fd_sc_hd__or2_4 _3730_ (.A(_3442_),
    .B(_3497_),
    .X(_3528_));
 sky130_fd_sc_hd__or3_1 _3731_ (.A(\as1802.instr_latch[5] ),
    .B(net163),
    .C(_3523_),
    .X(_3529_));
 sky130_fd_sc_hd__and3_1 _3732_ (.A(_3526_),
    .B(_3528_),
    .C(_3529_),
    .X(_3530_));
 sky130_fd_sc_hd__or3_1 _3733_ (.A(net827),
    .B(net809),
    .C(net852),
    .X(_3531_));
 sky130_fd_sc_hd__nand2_1 _3734_ (.A(_3499_),
    .B(_3531_),
    .Y(_3532_));
 sky130_fd_sc_hd__nor2_1 _3735_ (.A(net102),
    .B(_3532_),
    .Y(_3533_));
 sky130_fd_sc_hd__and3_1 _3736_ (.A(net209),
    .B(_3530_),
    .C(_3533_),
    .X(_3534_));
 sky130_fd_sc_hd__a32o_1 _3737_ (.A1(\as1802.instr_cycle[1] ),
    .A2(_3521_),
    .A3(_3534_),
    .B1(net274),
    .B2(_3491_),
    .X(_0015_));
 sky130_fd_sc_hd__and2b_2 _3738_ (.A_N(net39),
    .B(net46),
    .X(_3535_));
 sky130_fd_sc_hd__nor2_1 _3739_ (.A(net67),
    .B(_3535_),
    .Y(_3536_));
 sky130_fd_sc_hd__nor2_2 _3740_ (.A(_3432_),
    .B(net830),
    .Y(_3537_));
 sky130_fd_sc_hd__and2b_1 _3741_ (.A_N(_3536_),
    .B(_3537_),
    .X(_3538_));
 sky130_fd_sc_hd__or3_2 _3742_ (.A(_3432_),
    .B(\as1802.will_interrupt ),
    .C(_3536_),
    .X(_3539_));
 sky130_fd_sc_hd__nand2_2 _3743_ (.A(net173),
    .B(net830),
    .Y(_3540_));
 sky130_fd_sc_hd__nor2_2 _3744_ (.A(net833),
    .B(_3540_),
    .Y(_3541_));
 sky130_fd_sc_hd__o21a_1 _3745_ (.A1(_3538_),
    .A2(_3541_),
    .B1(net104),
    .X(_3542_));
 sky130_fd_sc_hd__nand2_2 _3746_ (.A(_3457_),
    .B(net352),
    .Y(_3543_));
 sky130_fd_sc_hd__or2_2 _3747_ (.A(_3456_),
    .B(_3543_),
    .X(_3544_));
 sky130_fd_sc_hd__nor3_1 _3748_ (.A(net171),
    .B(net366),
    .C(_3544_),
    .Y(_3545_));
 sky130_fd_sc_hd__nor2_1 _3749_ (.A(net356),
    .B(_3457_),
    .Y(_3546_));
 sky130_fd_sc_hd__and2_2 _3750_ (.A(_3456_),
    .B(net352),
    .X(_3547_));
 sky130_fd_sc_hd__nand2_4 _3751_ (.A(_3456_),
    .B(net352),
    .Y(_3548_));
 sky130_fd_sc_hd__nor2_1 _3752_ (.A(_3456_),
    .B(_3457_),
    .Y(_3549_));
 sky130_fd_sc_hd__nor2_8 _3753_ (.A(net356),
    .B(_3543_),
    .Y(_3550_));
 sky130_fd_sc_hd__or2_1 _3754_ (.A(net356),
    .B(_3543_),
    .X(_3551_));
 sky130_fd_sc_hd__nor2_2 _3755_ (.A(net172),
    .B(net102),
    .Y(_3552_));
 sky130_fd_sc_hd__nand2_4 _3756_ (.A(_3432_),
    .B(net105),
    .Y(_3553_));
 sky130_fd_sc_hd__or3_1 _3757_ (.A(_3549_),
    .B(_3550_),
    .C(_3552_),
    .X(_3554_));
 sky130_fd_sc_hd__nor2_1 _3758_ (.A(_3456_),
    .B(net352),
    .Y(_3555_));
 sky130_fd_sc_hd__nor2_1 _3759_ (.A(_3456_),
    .B(\as1802.mem_cycle[1] ),
    .Y(_3556_));
 sky130_fd_sc_hd__a221oi_4 _3760_ (.A1(_3457_),
    .A2(_3555_),
    .B1(_3556_),
    .B2(net366),
    .C1(_3546_),
    .Y(_3557_));
 sky130_fd_sc_hd__nand2_1 _3761_ (.A(net210),
    .B(_3557_),
    .Y(_3558_));
 sky130_fd_sc_hd__or4_2 _3762_ (.A(_3542_),
    .B(_3545_),
    .C(_3554_),
    .D(_3558_),
    .X(_3559_));
 sky130_fd_sc_hd__or3_1 _3763_ (.A(net830),
    .B(net103),
    .C(_3559_),
    .X(_3560_));
 sky130_fd_sc_hd__a21bo_1 _3764_ (.A1(net171),
    .A2(_3491_),
    .B1_N(_3560_),
    .X(_0014_));
 sky130_fd_sc_hd__nor2_2 _3765_ (.A(net164),
    .B(net167),
    .Y(_3561_));
 sky130_fd_sc_hd__or2_1 _3766_ (.A(net166),
    .B(\as1802.instr_latch[2] ),
    .X(_3562_));
 sky130_fd_sc_hd__and2_2 _3767_ (.A(net164),
    .B(net167),
    .X(_3563_));
 sky130_fd_sc_hd__or4_1 _3768_ (.A(net130),
    .B(net132),
    .C(net133),
    .D(net135),
    .X(_3564_));
 sky130_fd_sc_hd__or4_1 _3769_ (.A(net120),
    .B(net123),
    .C(net126),
    .D(net127),
    .X(_3565_));
 sky130_fd_sc_hd__or2_1 _3770_ (.A(_3564_),
    .B(_3565_),
    .X(_3566_));
 sky130_fd_sc_hd__nor3_1 _3771_ (.A(_3561_),
    .B(_3563_),
    .C(_3566_),
    .Y(_3567_));
 sky130_fd_sc_hd__o21a_1 _3772_ (.A1(_3561_),
    .A2(_3563_),
    .B1(_3566_),
    .X(_3568_));
 sky130_fd_sc_hd__or2_2 _3773_ (.A(net117),
    .B(net167),
    .X(_3569_));
 sky130_fd_sc_hd__nor2_4 _3774_ (.A(_3512_),
    .B(_3569_),
    .Y(_3570_));
 sky130_fd_sc_hd__inv_2 _3775_ (.A(_3570_),
    .Y(_3571_));
 sky130_fd_sc_hd__a21oi_1 _3776_ (.A1(net117),
    .A2(_3513_),
    .B1(_3570_),
    .Y(_3572_));
 sky130_fd_sc_hd__or2_1 _3777_ (.A(net63),
    .B(_3572_),
    .X(_3573_));
 sky130_fd_sc_hd__or4b_1 _3778_ (.A(net59),
    .B(_3561_),
    .C(_3563_),
    .D_N(_3508_),
    .X(_3574_));
 sky130_fd_sc_hd__a31o_1 _3779_ (.A1(net46),
    .A2(_3502_),
    .A3(_3563_),
    .B1(net161),
    .X(_3575_));
 sky130_fd_sc_hd__and2_2 _3780_ (.A(_3502_),
    .B(_3561_),
    .X(_3576_));
 sky130_fd_sc_hd__nor2_2 _3781_ (.A(net169),
    .B(_3569_),
    .Y(_3577_));
 sky130_fd_sc_hd__or2_2 _3782_ (.A(net169),
    .B(_3569_),
    .X(_3578_));
 sky130_fd_sc_hd__nor2_4 _3783_ (.A(net315),
    .B(_3578_),
    .Y(_3579_));
 sky130_fd_sc_hd__or2_2 _3784_ (.A(_3576_),
    .B(_3579_),
    .X(_3580_));
 sky130_fd_sc_hd__a22o_1 _3785_ (.A1(net59),
    .A2(_3508_),
    .B1(_3511_),
    .B2(net63),
    .X(_3581_));
 sky130_fd_sc_hd__o21ai_1 _3786_ (.A1(_3561_),
    .A2(_3563_),
    .B1(_3581_),
    .Y(_3582_));
 sky130_fd_sc_hd__and4bb_1 _3787_ (.A_N(_3575_),
    .B_N(_3580_),
    .C(_3582_),
    .D(_3574_),
    .X(_3583_));
 sky130_fd_sc_hd__o311a_2 _3788_ (.A1(_3516_),
    .A2(_3567_),
    .A3(_3568_),
    .B1(_3573_),
    .C1(_3583_),
    .X(_3584_));
 sky130_fd_sc_hd__mux4_1 _3789_ (.A0(\as1802.regs[8][14] ),
    .A1(\as1802.regs[9][14] ),
    .A2(\as1802.regs[10][14] ),
    .A3(\as1802.regs[11][14] ),
    .S0(net192),
    .S1(net188),
    .X(_3585_));
 sky130_fd_sc_hd__mux4_1 _3790_ (.A0(\as1802.regs[12][14] ),
    .A1(\as1802.regs[13][14] ),
    .A2(\as1802.regs[14][14] ),
    .A3(\as1802.regs[15][14] ),
    .S0(net192),
    .S1(net188),
    .X(_3586_));
 sky130_fd_sc_hd__nor2_1 _3791_ (.A(net115),
    .B(_3586_),
    .Y(_3587_));
 sky130_fd_sc_hd__mux4_1 _3792_ (.A0(\as1802.regs[4][14] ),
    .A1(\as1802.regs[5][14] ),
    .A2(\as1802.regs[6][14] ),
    .A3(\as1802.regs[7][14] ),
    .S0(net193),
    .S1(net189),
    .X(_3588_));
 sky130_fd_sc_hd__mux4_1 _3793_ (.A0(\as1802.regs[0][14] ),
    .A1(\as1802.regs[1][14] ),
    .A2(\as1802.regs[2][14] ),
    .A3(\as1802.regs[3][14] ),
    .S0(net193),
    .S1(net189),
    .X(_3589_));
 sky130_fd_sc_hd__mux2_1 _3794_ (.A0(_3588_),
    .A1(_3589_),
    .S(net115),
    .X(_3590_));
 sky130_fd_sc_hd__o21ai_1 _3795_ (.A1(net185),
    .A2(_3585_),
    .B1(_0003_),
    .Y(_3591_));
 sky130_fd_sc_hd__o2bb2a_4 _3796_ (.A1_N(net114),
    .A2_N(_3590_),
    .B1(_3591_),
    .B2(_3587_),
    .X(_3592_));
 sky130_fd_sc_hd__mux4_1 _3797_ (.A0(\as1802.regs[8][13] ),
    .A1(\as1802.regs[9][13] ),
    .A2(\as1802.regs[10][13] ),
    .A3(\as1802.regs[11][13] ),
    .S0(net192),
    .S1(net188),
    .X(_3593_));
 sky130_fd_sc_hd__nand2_1 _3798_ (.A(net116),
    .B(_3593_),
    .Y(_3594_));
 sky130_fd_sc_hd__mux4_1 _3799_ (.A0(\as1802.regs[12][13] ),
    .A1(\as1802.regs[13][13] ),
    .A2(\as1802.regs[14][13] ),
    .A3(\as1802.regs[15][13] ),
    .S0(net192),
    .S1(net188),
    .X(_3595_));
 sky130_fd_sc_hd__mux4_1 _3800_ (.A0(\as1802.regs[4][13] ),
    .A1(\as1802.regs[5][13] ),
    .A2(\as1802.regs[6][13] ),
    .A3(\as1802.regs[7][13] ),
    .S0(net192),
    .S1(net188),
    .X(_3596_));
 sky130_fd_sc_hd__mux4_1 _3801_ (.A0(\as1802.regs[0][13] ),
    .A1(\as1802.regs[1][13] ),
    .A2(\as1802.regs[2][13] ),
    .A3(\as1802.regs[3][13] ),
    .S0(net193),
    .S1(net189),
    .X(_3597_));
 sky130_fd_sc_hd__mux2_1 _3802_ (.A0(_3596_),
    .A1(_3597_),
    .S(net116),
    .X(_3598_));
 sky130_fd_sc_hd__a21oi_1 _3803_ (.A1(net185),
    .A2(_3595_),
    .B1(net114),
    .Y(_3599_));
 sky130_fd_sc_hd__a2bb2o_4 _3804_ (.A1_N(_0003_),
    .A2_N(_3598_),
    .B1(_3599_),
    .B2(_3594_),
    .X(_3600_));
 sky130_fd_sc_hd__mux4_1 _3805_ (.A0(\as1802.regs[8][12] ),
    .A1(\as1802.regs[9][12] ),
    .A2(\as1802.regs[10][12] ),
    .A3(\as1802.regs[11][12] ),
    .S0(net192),
    .S1(net188),
    .X(_3601_));
 sky130_fd_sc_hd__nand2_1 _3806_ (.A(net116),
    .B(_3601_),
    .Y(_3602_));
 sky130_fd_sc_hd__mux4_1 _3807_ (.A0(\as1802.regs[12][12] ),
    .A1(\as1802.regs[13][12] ),
    .A2(\as1802.regs[14][12] ),
    .A3(\as1802.regs[15][12] ),
    .S0(net192),
    .S1(net188),
    .X(_3603_));
 sky130_fd_sc_hd__mux4_1 _3808_ (.A0(\as1802.regs[4][12] ),
    .A1(\as1802.regs[5][12] ),
    .A2(\as1802.regs[6][12] ),
    .A3(\as1802.regs[7][12] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_3604_));
 sky130_fd_sc_hd__mux4_1 _3809_ (.A0(\as1802.regs[0][12] ),
    .A1(\as1802.regs[1][12] ),
    .A2(\as1802.regs[2][12] ),
    .A3(\as1802.regs[3][12] ),
    .S0(net193),
    .S1(net189),
    .X(_3605_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(_3604_),
    .A1(_3605_),
    .S(net116),
    .X(_3606_));
 sky130_fd_sc_hd__a21oi_1 _3811_ (.A1(net185),
    .A2(_3603_),
    .B1(net114),
    .Y(_3607_));
 sky130_fd_sc_hd__a2bb2o_4 _3812_ (.A1_N(_0003_),
    .A2_N(_3606_),
    .B1(_3607_),
    .B2(_3602_),
    .X(_3608_));
 sky130_fd_sc_hd__mux4_1 _3813_ (.A0(\as1802.regs[8][9] ),
    .A1(\as1802.regs[9][9] ),
    .A2(\as1802.regs[10][9] ),
    .A3(\as1802.regs[11][9] ),
    .S0(net192),
    .S1(net188),
    .X(_3609_));
 sky130_fd_sc_hd__nand2_1 _3814_ (.A(net116),
    .B(_3609_),
    .Y(_3610_));
 sky130_fd_sc_hd__mux4_1 _3815_ (.A0(\as1802.regs[12][9] ),
    .A1(\as1802.regs[13][9] ),
    .A2(\as1802.regs[14][9] ),
    .A3(\as1802.regs[15][9] ),
    .S0(net192),
    .S1(net188),
    .X(_3611_));
 sky130_fd_sc_hd__mux4_1 _3816_ (.A0(\as1802.regs[4][9] ),
    .A1(\as1802.regs[5][9] ),
    .A2(\as1802.regs[6][9] ),
    .A3(\as1802.regs[7][9] ),
    .S0(net192),
    .S1(net188),
    .X(_3612_));
 sky130_fd_sc_hd__mux4_1 _3817_ (.A0(\as1802.regs[0][9] ),
    .A1(\as1802.regs[1][9] ),
    .A2(\as1802.regs[2][9] ),
    .A3(\as1802.regs[3][9] ),
    .S0(net193),
    .S1(net189),
    .X(_3613_));
 sky130_fd_sc_hd__mux2_1 _3818_ (.A0(_3612_),
    .A1(_3613_),
    .S(net115),
    .X(_3614_));
 sky130_fd_sc_hd__a21oi_1 _3819_ (.A1(net185),
    .A2(_3611_),
    .B1(net114),
    .Y(_3615_));
 sky130_fd_sc_hd__a2bb2o_4 _3820_ (.A1_N(_0003_),
    .A2_N(_3614_),
    .B1(_3615_),
    .B2(_3610_),
    .X(_3616_));
 sky130_fd_sc_hd__mux4_1 _3821_ (.A0(\as1802.regs[8][8] ),
    .A1(\as1802.regs[9][8] ),
    .A2(\as1802.regs[10][8] ),
    .A3(\as1802.regs[11][8] ),
    .S0(net192),
    .S1(net188),
    .X(_3617_));
 sky130_fd_sc_hd__mux4_1 _3822_ (.A0(\as1802.regs[12][8] ),
    .A1(\as1802.regs[13][8] ),
    .A2(\as1802.regs[14][8] ),
    .A3(\as1802.regs[15][8] ),
    .S0(net192),
    .S1(net188),
    .X(_3618_));
 sky130_fd_sc_hd__mux2_1 _3823_ (.A0(_3617_),
    .A1(_3618_),
    .S(net185),
    .X(_3619_));
 sky130_fd_sc_hd__mux4_1 _3824_ (.A0(\as1802.regs[4][8] ),
    .A1(\as1802.regs[5][8] ),
    .A2(\as1802.regs[6][8] ),
    .A3(\as1802.regs[7][8] ),
    .S0(net193),
    .S1(net189),
    .X(_3620_));
 sky130_fd_sc_hd__mux4_1 _3825_ (.A0(\as1802.regs[0][8] ),
    .A1(\as1802.regs[1][8] ),
    .A2(\as1802.regs[2][8] ),
    .A3(\as1802.regs[3][8] ),
    .S0(net193),
    .S1(net189),
    .X(_3621_));
 sky130_fd_sc_hd__mux2_1 _3826_ (.A0(_3620_),
    .A1(_3621_),
    .S(net116),
    .X(_3622_));
 sky130_fd_sc_hd__mux2_4 _3827_ (.A0(_3619_),
    .A1(_3622_),
    .S(net114),
    .X(_3623_));
 sky130_fd_sc_hd__mux4_1 _3828_ (.A0(\as1802.regs[8][5] ),
    .A1(\as1802.regs[9][5] ),
    .A2(\as1802.regs[10][5] ),
    .A3(\as1802.regs[11][5] ),
    .S0(net191),
    .S1(net187),
    .X(_3624_));
 sky130_fd_sc_hd__nand2_1 _3829_ (.A(net115),
    .B(_3624_),
    .Y(_3625_));
 sky130_fd_sc_hd__mux4_1 _3830_ (.A0(\as1802.regs[12][5] ),
    .A1(\as1802.regs[13][5] ),
    .A2(\as1802.regs[14][5] ),
    .A3(\as1802.regs[15][5] ),
    .S0(net190),
    .S1(net186),
    .X(_3626_));
 sky130_fd_sc_hd__mux4_1 _3831_ (.A0(\as1802.regs[4][5] ),
    .A1(\as1802.regs[5][5] ),
    .A2(\as1802.regs[6][5] ),
    .A3(\as1802.regs[7][5] ),
    .S0(net190),
    .S1(net186),
    .X(_3627_));
 sky130_fd_sc_hd__mux4_1 _3832_ (.A0(\as1802.regs[0][5] ),
    .A1(\as1802.regs[1][5] ),
    .A2(\as1802.regs[2][5] ),
    .A3(\as1802.regs[3][5] ),
    .S0(net191),
    .S1(net187),
    .X(_3628_));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(_3627_),
    .A1(_3628_),
    .S(net115),
    .X(_3629_));
 sky130_fd_sc_hd__a21oi_1 _3834_ (.A1(net185),
    .A2(_3626_),
    .B1(net114),
    .Y(_0387_));
 sky130_fd_sc_hd__a2bb2o_2 _3835_ (.A1_N(_0003_),
    .A2_N(_3629_),
    .B1(_0387_),
    .B2(_3625_),
    .X(_0388_));
 sky130_fd_sc_hd__mux4_1 _3836_ (.A0(\as1802.regs[8][4] ),
    .A1(\as1802.regs[9][4] ),
    .A2(\as1802.regs[10][4] ),
    .A3(\as1802.regs[11][4] ),
    .S0(net190),
    .S1(net186),
    .X(_0389_));
 sky130_fd_sc_hd__mux4_1 _3837_ (.A0(\as1802.regs[12][4] ),
    .A1(\as1802.regs[13][4] ),
    .A2(\as1802.regs[14][4] ),
    .A3(\as1802.regs[15][4] ),
    .S0(net190),
    .S1(net186),
    .X(_0390_));
 sky130_fd_sc_hd__nor2_1 _3838_ (.A(net115),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__mux4_1 _3839_ (.A0(\as1802.regs[4][4] ),
    .A1(\as1802.regs[5][4] ),
    .A2(\as1802.regs[6][4] ),
    .A3(\as1802.regs[7][4] ),
    .S0(net190),
    .S1(net186),
    .X(_0392_));
 sky130_fd_sc_hd__mux4_1 _3840_ (.A0(\as1802.regs[0][4] ),
    .A1(\as1802.regs[1][4] ),
    .A2(\as1802.regs[2][4] ),
    .A3(\as1802.regs[3][4] ),
    .S0(net191),
    .S1(net187),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3841_ (.A0(_0392_),
    .A1(_0393_),
    .S(net115),
    .X(_0394_));
 sky130_fd_sc_hd__o21ai_1 _3842_ (.A1(net185),
    .A2(_0389_),
    .B1(_0003_),
    .Y(_0395_));
 sky130_fd_sc_hd__o2bb2a_2 _3843_ (.A1_N(net114),
    .A2_N(_0394_),
    .B1(_0395_),
    .B2(_0391_),
    .X(_0396_));
 sky130_fd_sc_hd__mux4_1 _3844_ (.A0(\as1802.regs[8][3] ),
    .A1(\as1802.regs[9][3] ),
    .A2(\as1802.regs[10][3] ),
    .A3(\as1802.regs[11][3] ),
    .S0(net190),
    .S1(net186),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _3845_ (.A(net115),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__mux4_1 _3846_ (.A0(\as1802.regs[12][3] ),
    .A1(\as1802.regs[13][3] ),
    .A2(\as1802.regs[14][3] ),
    .A3(\as1802.regs[15][3] ),
    .S0(net190),
    .S1(net186),
    .X(_0399_));
 sky130_fd_sc_hd__mux4_1 _3847_ (.A0(\as1802.regs[4][3] ),
    .A1(\as1802.regs[5][3] ),
    .A2(\as1802.regs[6][3] ),
    .A3(\as1802.regs[7][3] ),
    .S0(net190),
    .S1(net186),
    .X(_0400_));
 sky130_fd_sc_hd__mux4_1 _3848_ (.A0(\as1802.regs[0][3] ),
    .A1(\as1802.regs[1][3] ),
    .A2(\as1802.regs[2][3] ),
    .A3(\as1802.regs[3][3] ),
    .S0(net191),
    .S1(net187),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3849_ (.A0(_0400_),
    .A1(_0401_),
    .S(net115),
    .X(_0402_));
 sky130_fd_sc_hd__a21oi_1 _3850_ (.A1(net185),
    .A2(_0399_),
    .B1(net114),
    .Y(_0403_));
 sky130_fd_sc_hd__a2bb2o_2 _3851_ (.A1_N(_0003_),
    .A2_N(_0402_),
    .B1(_0403_),
    .B2(_0398_),
    .X(_0404_));
 sky130_fd_sc_hd__mux4_1 _3852_ (.A0(\as1802.regs[8][2] ),
    .A1(\as1802.regs[9][2] ),
    .A2(\as1802.regs[10][2] ),
    .A3(\as1802.regs[11][2] ),
    .S0(net190),
    .S1(net186),
    .X(_0405_));
 sky130_fd_sc_hd__mux4_1 _3853_ (.A0(\as1802.regs[12][2] ),
    .A1(\as1802.regs[13][2] ),
    .A2(\as1802.regs[14][2] ),
    .A3(\as1802.regs[15][2] ),
    .S0(net190),
    .S1(net186),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _3854_ (.A(net115),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _3855_ (.A0(\as1802.regs[4][2] ),
    .A1(\as1802.regs[5][2] ),
    .A2(\as1802.regs[6][2] ),
    .A3(\as1802.regs[7][2] ),
    .S0(net191),
    .S1(net187),
    .X(_0408_));
 sky130_fd_sc_hd__mux4_1 _3856_ (.A0(\as1802.regs[0][2] ),
    .A1(\as1802.regs[1][2] ),
    .A2(\as1802.regs[2][2] ),
    .A3(\as1802.regs[3][2] ),
    .S0(net191),
    .S1(net187),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3857_ (.A0(_0408_),
    .A1(_0409_),
    .S(net115),
    .X(_0410_));
 sky130_fd_sc_hd__o211a_1 _3858_ (.A1(net185),
    .A2(_0405_),
    .B1(_0407_),
    .C1(_0003_),
    .X(_0411_));
 sky130_fd_sc_hd__a21oi_4 _3859_ (.A1(net114),
    .A2(_0410_),
    .B1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__mux4_1 _3860_ (.A0(\as1802.regs[8][0] ),
    .A1(\as1802.regs[9][0] ),
    .A2(\as1802.regs[10][0] ),
    .A3(\as1802.regs[11][0] ),
    .S0(net190),
    .S1(net186),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _3861_ (.A(net185),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__mux4_1 _3862_ (.A0(\as1802.regs[12][0] ),
    .A1(\as1802.regs[13][0] ),
    .A2(\as1802.regs[14][0] ),
    .A3(\as1802.regs[15][0] ),
    .S0(net190),
    .S1(net186),
    .X(_0415_));
 sky130_fd_sc_hd__mux4_1 _3863_ (.A0(\as1802.regs[4][0] ),
    .A1(\as1802.regs[5][0] ),
    .A2(\as1802.regs[6][0] ),
    .A3(\as1802.regs[7][0] ),
    .S0(net191),
    .S1(net187),
    .X(_0416_));
 sky130_fd_sc_hd__mux4_1 _3864_ (.A0(\as1802.regs[0][0] ),
    .A1(\as1802.regs[1][0] ),
    .A2(\as1802.regs[2][0] ),
    .A3(\as1802.regs[3][0] ),
    .S0(net191),
    .S1(net187),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(_0416_),
    .A1(_0417_),
    .S(net115),
    .X(_0418_));
 sky130_fd_sc_hd__o21ai_1 _3866_ (.A1(net115),
    .A2(_0415_),
    .B1(_0003_),
    .Y(_0419_));
 sky130_fd_sc_hd__o2bb2a_4 _3867_ (.A1_N(net114),
    .A2_N(_0418_),
    .B1(_0419_),
    .B2(_0414_),
    .X(_0420_));
 sky130_fd_sc_hd__mux4_1 _3868_ (.A0(\as1802.regs[8][1] ),
    .A1(\as1802.regs[9][1] ),
    .A2(\as1802.regs[10][1] ),
    .A3(\as1802.regs[11][1] ),
    .S0(net190),
    .S1(net186),
    .X(_0421_));
 sky130_fd_sc_hd__mux4_1 _3869_ (.A0(\as1802.regs[12][1] ),
    .A1(\as1802.regs[13][1] ),
    .A2(\as1802.regs[14][1] ),
    .A3(\as1802.regs[15][1] ),
    .S0(net190),
    .S1(net186),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3870_ (.A0(_0421_),
    .A1(_0422_),
    .S(net185),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _3871_ (.A(_0003_),
    .B(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__mux4_1 _3872_ (.A0(\as1802.regs[4][1] ),
    .A1(\as1802.regs[5][1] ),
    .A2(\as1802.regs[6][1] ),
    .A3(\as1802.regs[7][1] ),
    .S0(net191),
    .S1(net187),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_1 _3873_ (.A0(\as1802.regs[0][1] ),
    .A1(\as1802.regs[1][1] ),
    .A2(\as1802.regs[2][1] ),
    .A3(\as1802.regs[3][1] ),
    .S0(net191),
    .S1(net187),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(_0425_),
    .A1(_0426_),
    .S(net115),
    .X(_0427_));
 sky130_fd_sc_hd__a21oi_4 _3875_ (.A1(net114),
    .A2(_0427_),
    .B1(_0424_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_0420_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__and3_1 _3877_ (.A(_0412_),
    .B(_0420_),
    .C(_0428_),
    .X(_0430_));
 sky130_fd_sc_hd__and2_1 _3878_ (.A(_0404_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__and3_1 _3879_ (.A(_0396_),
    .B(_0404_),
    .C(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__and2_1 _3880_ (.A(_0388_),
    .B(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__mux4_1 _3881_ (.A0(\as1802.regs[8][6] ),
    .A1(\as1802.regs[9][6] ),
    .A2(\as1802.regs[10][6] ),
    .A3(\as1802.regs[11][6] ),
    .S0(net190),
    .S1(net186),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_1 _3882_ (.A(net185),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__mux4_1 _3883_ (.A0(\as1802.regs[12][6] ),
    .A1(\as1802.regs[13][6] ),
    .A2(\as1802.regs[14][6] ),
    .A3(\as1802.regs[15][6] ),
    .S0(net190),
    .S1(net186),
    .X(_0436_));
 sky130_fd_sc_hd__mux4_1 _3884_ (.A0(\as1802.regs[4][6] ),
    .A1(\as1802.regs[5][6] ),
    .A2(\as1802.regs[6][6] ),
    .A3(\as1802.regs[7][6] ),
    .S0(net191),
    .S1(net187),
    .X(_0437_));
 sky130_fd_sc_hd__mux4_1 _3885_ (.A0(\as1802.regs[0][6] ),
    .A1(\as1802.regs[1][6] ),
    .A2(\as1802.regs[2][6] ),
    .A3(\as1802.regs[3][6] ),
    .S0(net191),
    .S1(net187),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3886_ (.A0(_0437_),
    .A1(_0438_),
    .S(net115),
    .X(_0439_));
 sky130_fd_sc_hd__o21ai_1 _3887_ (.A1(net115),
    .A2(_0436_),
    .B1(_0003_),
    .Y(_0440_));
 sky130_fd_sc_hd__o2bb2a_4 _3888_ (.A1_N(net114),
    .A2_N(_0439_),
    .B1(_0440_),
    .B2(_0435_),
    .X(_0441_));
 sky130_fd_sc_hd__inv_2 _3889_ (.A(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__and3_1 _3890_ (.A(_0388_),
    .B(_0432_),
    .C(_0441_),
    .X(_0443_));
 sky130_fd_sc_hd__mux4_1 _3891_ (.A0(\as1802.regs[8][7] ),
    .A1(\as1802.regs[9][7] ),
    .A2(\as1802.regs[10][7] ),
    .A3(\as1802.regs[11][7] ),
    .S0(net191),
    .S1(net187),
    .X(_0444_));
 sky130_fd_sc_hd__mux4_1 _3892_ (.A0(\as1802.regs[12][7] ),
    .A1(\as1802.regs[13][7] ),
    .A2(\as1802.regs[14][7] ),
    .A3(\as1802.regs[15][7] ),
    .S0(net191),
    .S1(net187),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3893_ (.A0(_0444_),
    .A1(_0445_),
    .S(net185),
    .X(_0446_));
 sky130_fd_sc_hd__and2_1 _3894_ (.A(_0003_),
    .B(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__mux4_1 _3895_ (.A0(\as1802.regs[4][7] ),
    .A1(\as1802.regs[5][7] ),
    .A2(\as1802.regs[6][7] ),
    .A3(\as1802.regs[7][7] ),
    .S0(_0000_),
    .S1(_0001_),
    .X(_0448_));
 sky130_fd_sc_hd__mux4_1 _3896_ (.A0(\as1802.regs[0][7] ),
    .A1(\as1802.regs[1][7] ),
    .A2(\as1802.regs[2][7] ),
    .A3(\as1802.regs[3][7] ),
    .S0(net191),
    .S1(net187),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(_0448_),
    .A1(_0449_),
    .S(net116),
    .X(_0450_));
 sky130_fd_sc_hd__a21oi_4 _3898_ (.A1(_3467_),
    .A2(_0450_),
    .B1(_0447_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _3899_ (.A(_0443_),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _3900_ (.A(_3623_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__and2_1 _3901_ (.A(_3616_),
    .B(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__mux4_1 _3902_ (.A0(\as1802.regs[8][10] ),
    .A1(\as1802.regs[9][10] ),
    .A2(\as1802.regs[10][10] ),
    .A3(\as1802.regs[11][10] ),
    .S0(net192),
    .S1(net188),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _3903_ (.A(net185),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__mux4_1 _3904_ (.A0(\as1802.regs[12][10] ),
    .A1(\as1802.regs[13][10] ),
    .A2(\as1802.regs[14][10] ),
    .A3(\as1802.regs[15][10] ),
    .S0(net192),
    .S1(net188),
    .X(_0457_));
 sky130_fd_sc_hd__mux4_1 _3905_ (.A0(\as1802.regs[4][10] ),
    .A1(\as1802.regs[5][10] ),
    .A2(\as1802.regs[6][10] ),
    .A3(\as1802.regs[7][10] ),
    .S0(net192),
    .S1(net188),
    .X(_0458_));
 sky130_fd_sc_hd__mux4_1 _3906_ (.A0(\as1802.regs[0][10] ),
    .A1(\as1802.regs[1][10] ),
    .A2(\as1802.regs[2][10] ),
    .A3(\as1802.regs[3][10] ),
    .S0(net193),
    .S1(net189),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(_0458_),
    .A1(_0459_),
    .S(net116),
    .X(_0460_));
 sky130_fd_sc_hd__o21ai_1 _3908_ (.A1(net116),
    .A2(_0457_),
    .B1(_0003_),
    .Y(_0461_));
 sky130_fd_sc_hd__o2bb2a_4 _3909_ (.A1_N(net114),
    .A2_N(_0460_),
    .B1(_0461_),
    .B2(_0456_),
    .X(_0462_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_0454_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__mux4_1 _3911_ (.A0(\as1802.regs[8][11] ),
    .A1(\as1802.regs[9][11] ),
    .A2(\as1802.regs[10][11] ),
    .A3(\as1802.regs[11][11] ),
    .S0(net193),
    .S1(net189),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _3912_ (.A(net116),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__mux4_1 _3913_ (.A0(\as1802.regs[12][11] ),
    .A1(\as1802.regs[13][11] ),
    .A2(\as1802.regs[14][11] ),
    .A3(\as1802.regs[15][11] ),
    .S0(net192),
    .S1(net188),
    .X(_0466_));
 sky130_fd_sc_hd__mux4_1 _3914_ (.A0(\as1802.regs[4][11] ),
    .A1(\as1802.regs[5][11] ),
    .A2(\as1802.regs[6][11] ),
    .A3(\as1802.regs[7][11] ),
    .S0(net193),
    .S1(net189),
    .X(_0467_));
 sky130_fd_sc_hd__and2_1 _3915_ (.A(net185),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__mux4_1 _3916_ (.A0(\as1802.regs[0][11] ),
    .A1(\as1802.regs[1][11] ),
    .A2(\as1802.regs[2][11] ),
    .A3(\as1802.regs[3][11] ),
    .S0(net193),
    .S1(net189),
    .X(_0469_));
 sky130_fd_sc_hd__a21oi_1 _3917_ (.A1(net116),
    .A2(_0469_),
    .B1(_0468_),
    .Y(_0470_));
 sky130_fd_sc_hd__a21o_1 _3918_ (.A1(_0002_),
    .A2(_0466_),
    .B1(net114),
    .X(_0471_));
 sky130_fd_sc_hd__a2bb2o_2 _3919_ (.A1_N(_0471_),
    .A2_N(_0465_),
    .B1(net114),
    .B2(_0470_),
    .X(_0472_));
 sky130_fd_sc_hd__o2bb2a_2 _3920_ (.A1_N(_3467_),
    .A2_N(_0470_),
    .B1(_0471_),
    .B2(_0465_),
    .X(_0473_));
 sky130_fd_sc_hd__nor2_1 _3921_ (.A(_0463_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__and2_1 _3922_ (.A(_3608_),
    .B(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__and3_1 _3923_ (.A(_3600_),
    .B(_3608_),
    .C(_0474_),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _3924_ (.A(_3592_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__mux4_1 _3925_ (.A0(\as1802.regs[8][15] ),
    .A1(\as1802.regs[9][15] ),
    .A2(\as1802.regs[10][15] ),
    .A3(\as1802.regs[11][15] ),
    .S0(net193),
    .S1(net189),
    .X(_0478_));
 sky130_fd_sc_hd__mux4_1 _3926_ (.A0(\as1802.regs[12][15] ),
    .A1(\as1802.regs[13][15] ),
    .A2(\as1802.regs[14][15] ),
    .A3(\as1802.regs[15][15] ),
    .S0(net193),
    .S1(net189),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(_0478_),
    .A1(_0479_),
    .S(_0002_),
    .X(_0480_));
 sky130_fd_sc_hd__and2_1 _3928_ (.A(_0003_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__mux4_1 _3929_ (.A0(\as1802.regs[4][15] ),
    .A1(\as1802.regs[5][15] ),
    .A2(\as1802.regs[6][15] ),
    .A3(\as1802.regs[7][15] ),
    .S0(net193),
    .S1(net189),
    .X(_0482_));
 sky130_fd_sc_hd__mux4_1 _3930_ (.A0(\as1802.regs[0][15] ),
    .A1(\as1802.regs[1][15] ),
    .A2(\as1802.regs[2][15] ),
    .A3(\as1802.regs[3][15] ),
    .S0(net193),
    .S1(net189),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(_0482_),
    .A1(_0483_),
    .S(net116),
    .X(_0484_));
 sky130_fd_sc_hd__a21oi_4 _3932_ (.A1(net114),
    .A2(_0484_),
    .B1(_0481_),
    .Y(_0485_));
 sky130_fd_sc_hd__xnor2_2 _3933_ (.A(_0477_),
    .B(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__or2_1 _3934_ (.A(_0454_),
    .B(_0462_),
    .X(_0487_));
 sky130_fd_sc_hd__and2_1 _3935_ (.A(_0463_),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__or2_1 _3936_ (.A(_0443_),
    .B(_0451_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _3937_ (.A(_0452_),
    .B(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(_0433_),
    .B(_0441_),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _3939_ (.A(_0443_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and4b_1 _3940_ (.A_N(_0420_),
    .B(_0428_),
    .C(_0396_),
    .D(_0412_),
    .X(_0493_));
 sky130_fd_sc_hd__and3_1 _3941_ (.A(net161),
    .B(_0404_),
    .C(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and4b_1 _3942_ (.A_N(_3623_),
    .B(_3592_),
    .C(_3616_),
    .D(_0388_),
    .X(_0495_));
 sky130_fd_sc_hd__and4_1 _3943_ (.A(_3600_),
    .B(_3608_),
    .C(_0472_),
    .D(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__and4bb_1 _3944_ (.A_N(_0490_),
    .B_N(_0492_),
    .C(_0494_),
    .D(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__a31oi_4 _3945_ (.A1(_0486_),
    .A2(_0488_),
    .A3(_0497_),
    .B1(_3584_),
    .Y(_0498_));
 sky130_fd_sc_hd__nor2_1 _3946_ (.A(net168),
    .B(_3516_),
    .Y(_0499_));
 sky130_fd_sc_hd__or2_4 _3947_ (.A(net167),
    .B(_3516_),
    .X(_0500_));
 sky130_fd_sc_hd__nor2_1 _3948_ (.A(_3566_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_4 _3949_ (.A(net167),
    .B(_3512_),
    .Y(_0502_));
 sky130_fd_sc_hd__a22o_1 _3950_ (.A1(\as1802.EF_l[0] ),
    .A2(_3503_),
    .B1(_0502_),
    .B2(net63),
    .X(_0503_));
 sky130_fd_sc_hd__a21o_1 _3951_ (.A1(\as1802.EF_l[2] ),
    .A2(_3517_),
    .B1(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _3952_ (.A1(\as1802.EF_l[1] ),
    .A2(net97),
    .B1(_3513_),
    .B2(\as1802.EF_l[3] ),
    .X(_0505_));
 sky130_fd_sc_hd__a211o_1 _3953_ (.A1(\as1802.instr_latch[0] ),
    .A2(_3445_),
    .B1(net167),
    .C1(net169),
    .X(_0506_));
 sky130_fd_sc_hd__or4b_1 _3954_ (.A(_0501_),
    .B(_0504_),
    .C(_0505_),
    .D_N(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__xnor2_1 _3955_ (.A(net117),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _3956_ (.A(net211),
    .B(net104),
    .Y(_0509_));
 sky130_fd_sc_hd__and3_1 _3957_ (.A(\as1802.instr_latch[5] ),
    .B(\as1802.instr_latch[4] ),
    .C(_3494_),
    .X(_0510_));
 sky130_fd_sc_hd__and4bb_2 _3958_ (.A_N(_3517_),
    .B_N(_3580_),
    .C(_0510_),
    .D(net171),
    .X(_0511_));
 sky130_fd_sc_hd__and4_1 _3959_ (.A(_3440_),
    .B(\as1802.instr_latch[6] ),
    .C(\as1802.instr_latch[5] ),
    .D(net163),
    .X(_0512_));
 sky130_fd_sc_hd__or3_4 _3960_ (.A(_3441_),
    .B(_3442_),
    .C(_3523_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2b_1 _3961_ (.A_N(net167),
    .B(net169),
    .Y(_0514_));
 sky130_fd_sc_hd__and4_2 _3962_ (.A(net171),
    .B(_3516_),
    .C(_3569_),
    .D(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__and2_2 _3963_ (.A(net100),
    .B(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__or2_1 _3964_ (.A(_0511_),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__and4_1 _3965_ (.A(net210),
    .B(net104),
    .C(net96),
    .D(_0508_),
    .X(_0518_));
 sky130_fd_sc_hd__a31o_1 _3966_ (.A1(_3521_),
    .A2(_3534_),
    .A3(_0498_),
    .B1(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_1 _3967_ (.A1(net824),
    .A2(_3491_),
    .B1(_0519_),
    .B2(net171),
    .X(_0520_));
 sky130_fd_sc_hd__a31o_1 _3968_ (.A1(net210),
    .A2(net104),
    .A3(_0517_),
    .B1(_0520_),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _3969_ (.A(net171),
    .B(_3521_),
    .Y(_0521_));
 sky130_fd_sc_hd__and4b_1 _3970_ (.A_N(_0498_),
    .B(_3534_),
    .C(_3521_),
    .D(net732),
    .X(_0522_));
 sky130_fd_sc_hd__o21ai_1 _3971_ (.A1(_3463_),
    .A2(_3517_),
    .B1(_0510_),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_2 _3972_ (.A(_3580_),
    .B(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__nand2_1 _3973_ (.A(_3580_),
    .B(_0510_),
    .Y(_0525_));
 sky130_fd_sc_hd__nor2_2 _3974_ (.A(_0513_),
    .B(_0515_),
    .Y(_0526_));
 sky130_fd_sc_hd__or2_4 _3975_ (.A(_0513_),
    .B(_0515_),
    .X(_0527_));
 sky130_fd_sc_hd__nor2_2 _3976_ (.A(net161),
    .B(_3489_),
    .Y(_0528_));
 sky130_fd_sc_hd__o21a_1 _3977_ (.A1(\as1802.instr_cycle[1] ),
    .A2(net274),
    .B1(net96),
    .X(_0529_));
 sky130_fd_sc_hd__nand2_1 _3978_ (.A(_3442_),
    .B(_3485_),
    .Y(_0530_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(_3494_),
    .A1(_0530_),
    .S(\as1802.instr_latch[5] ),
    .X(_0531_));
 sky130_fd_sc_hd__and3_1 _3980_ (.A(_0524_),
    .B(_0525_),
    .C(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__or2_1 _3981_ (.A(_3442_),
    .B(_3531_),
    .X(_0533_));
 sky130_fd_sc_hd__or3_1 _3982_ (.A(_3441_),
    .B(net163),
    .C(_3495_),
    .X(_0534_));
 sky130_fd_sc_hd__nor2_4 _3983_ (.A(net852),
    .B(_3485_),
    .Y(_0535_));
 sky130_fd_sc_hd__nand2_4 _3984_ (.A(_3441_),
    .B(_3484_),
    .Y(_0536_));
 sky130_fd_sc_hd__or4b_1 _3985_ (.A(_0526_),
    .B(_0528_),
    .C(_0529_),
    .D_N(_0532_),
    .X(_0537_));
 sky130_fd_sc_hd__or2_1 _3986_ (.A(net163),
    .B(_3531_),
    .X(_0538_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(net104),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__and3_2 _3988_ (.A(_3499_),
    .B(_3529_),
    .C(_0533_),
    .X(_0540_));
 sky130_fd_sc_hd__and3b_1 _3989_ (.A_N(_0539_),
    .B(_0540_),
    .C(_3528_),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_2 _3990_ (.A(_3442_),
    .B(_3487_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(\as1802.instr_latch[4] ),
    .B(_3486_),
    .Y(_0543_));
 sky130_fd_sc_hd__or3_2 _3992_ (.A(\as1802.instr_latch[5] ),
    .B(_3442_),
    .C(_3495_),
    .X(_0544_));
 sky130_fd_sc_hd__nor2_1 _3993_ (.A(_0509_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a221o_1 _3994_ (.A1(net104),
    .A2(_0537_),
    .B1(_0541_),
    .B2(_0542_),
    .C1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__o31a_1 _3995_ (.A1(net732),
    .A2(\as1802.instr_cycle[1] ),
    .A3(net274),
    .B1(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__or3b_1 _3996_ (.A(\as1802.will_interrupt ),
    .B(net103),
    .C_N(_3536_),
    .X(_0548_));
 sky130_fd_sc_hd__a32o_1 _3997_ (.A1(net274),
    .A2(net104),
    .A3(_3496_),
    .B1(_0548_),
    .B2(net173),
    .X(_0549_));
 sky130_fd_sc_hd__nor2_2 _3998_ (.A(net171),
    .B(\as1802.instr_cycle[1] ),
    .Y(_0550_));
 sky130_fd_sc_hd__o221a_1 _3999_ (.A1(net732),
    .A2(\as1802.instr_cycle[1] ),
    .B1(_3506_),
    .B2(_3520_),
    .C1(_3501_),
    .X(_0551_));
 sky130_fd_sc_hd__a211o_1 _4000_ (.A1(_3534_),
    .A2(_0551_),
    .B1(_0549_),
    .C1(net206),
    .X(_0552_));
 sky130_fd_sc_hd__and4b_1 _4001_ (.A_N(_0508_),
    .B(net96),
    .C(net104),
    .D(net732),
    .X(_0553_));
 sky130_fd_sc_hd__or4_1 _4002_ (.A(_0522_),
    .B(net733),
    .C(_0552_),
    .D(_0553_),
    .X(_0012_));
 sky130_fd_sc_hd__a21o_2 _4003_ (.A1(net60),
    .A2(net19),
    .B1(\as1802.MRD ),
    .X(net56));
 sky130_fd_sc_hd__nor2_2 _4004_ (.A(clknet_leaf_12_wb_clk_i),
    .B(net17),
    .Y(_0554_));
 sky130_fd_sc_hd__a221o_2 _4005_ (.A1(net60),
    .A2(net20),
    .B1(net18),
    .B2(_0554_),
    .C1(net45),
    .X(_0555_));
 sky130_fd_sc_hd__a31o_2 _4006_ (.A1(clknet_leaf_12_wb_clk_i),
    .A2(net17),
    .A3(_3468_),
    .B1(_0555_),
    .X(net58));
 sky130_fd_sc_hd__or3_1 _4007_ (.A(_3485_),
    .B(_3492_),
    .C(_3553_),
    .X(_0556_));
 sky130_fd_sc_hd__or3_2 _4008_ (.A(net172),
    .B(net99),
    .C(_0535_),
    .X(_0557_));
 sky130_fd_sc_hd__nand2_1 _4009_ (.A(_3530_),
    .B(_3533_),
    .Y(_0558_));
 sky130_fd_sc_hd__nor2_1 _4010_ (.A(_0557_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__or2_1 _4011_ (.A(_0557_),
    .B(_0558_),
    .X(_0560_));
 sky130_fd_sc_hd__o211ai_1 _4012_ (.A1(_3440_),
    .A2(_3492_),
    .B1(_0559_),
    .C1(net809),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _4013_ (.A(_3488_),
    .B(_3552_),
    .Y(_0562_));
 sky130_fd_sc_hd__a21oi_1 _4014_ (.A1(_0556_),
    .A2(_0561_),
    .B1(net206),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(_3526_),
    .B(_0540_),
    .Y(_0564_));
 sky130_fd_sc_hd__o21ai_1 _4016_ (.A1(net102),
    .A2(_3528_),
    .B1(_0538_),
    .Y(_0565_));
 sky130_fd_sc_hd__a22o_1 _4017_ (.A1(_3552_),
    .A2(_0564_),
    .B1(_0565_),
    .B2(_3432_),
    .X(_0566_));
 sky130_fd_sc_hd__o41a_1 _4018_ (.A1(net102),
    .A2(_3537_),
    .A3(_3541_),
    .A4(_0566_),
    .B1(net209),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_4 _4019_ (.A(net172),
    .B(net206),
    .Y(_0568_));
 sky130_fd_sc_hd__nand2_4 _4020_ (.A(_3432_),
    .B(net211),
    .Y(_0569_));
 sky130_fd_sc_hd__nor2_8 _4021_ (.A(net102),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_4 _4022_ (.A(net104),
    .B(_0568_),
    .Y(_0571_));
 sky130_fd_sc_hd__and3_2 _4023_ (.A(net99),
    .B(_0515_),
    .C(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_4 _4024_ (.A(_0516_),
    .B(_0570_),
    .Y(_0573_));
 sky130_fd_sc_hd__nor2_4 _4025_ (.A(net163),
    .B(_0536_),
    .Y(_0574_));
 sky130_fd_sc_hd__and3_1 _4026_ (.A(_3432_),
    .B(_3442_),
    .C(_0535_),
    .X(_0575_));
 sky130_fd_sc_hd__inv_2 _4027_ (.A(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a31o_1 _4028_ (.A1(net211),
    .A2(_3533_),
    .A3(_0575_),
    .B1(_0572_),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_4 _4029_ (.A(_3442_),
    .B(_0536_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _4030_ (.A(net163),
    .B(_0535_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_1 _4031_ (.A(_3489_),
    .B(_0536_),
    .Y(_0580_));
 sky130_fd_sc_hd__or2_1 _4032_ (.A(net173),
    .B(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__or2_1 _4033_ (.A(_0544_),
    .B(_0557_),
    .X(_0582_));
 sky130_fd_sc_hd__nor2_1 _4034_ (.A(_3444_),
    .B(_3578_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_4 _4035_ (.A(net810),
    .B(_3577_),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_4 _4036_ (.A(net167),
    .B(net169),
    .Y(_0585_));
 sky130_fd_sc_hd__or2_4 _4037_ (.A(net168),
    .B(net170),
    .X(_0586_));
 sky130_fd_sc_hd__nand2_1 _4038_ (.A(net117),
    .B(_0585_),
    .Y(_0587_));
 sky130_fd_sc_hd__and4_1 _4039_ (.A(_3533_),
    .B(_0526_),
    .C(_0568_),
    .D(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__a2bb2o_1 _4040_ (.A1_N(_0509_),
    .A2_N(_0582_),
    .B1(_0584_),
    .B2(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__a31o_1 _4041_ (.A1(_3440_),
    .A2(\as1802.instr_latch[6] ),
    .A3(_3493_),
    .B1(net172),
    .X(_0590_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(_3440_),
    .B(_3553_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(_0534_),
    .B(_0544_),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2_1 _4044_ (.A(_3484_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a41o_1 _4045_ (.A1(net211),
    .A2(net95),
    .A3(_0591_),
    .A4(_0593_),
    .B1(_0563_),
    .X(_0594_));
 sky130_fd_sc_hd__or4_4 _4046_ (.A(_0567_),
    .B(_0577_),
    .C(_0589_),
    .D(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _4047_ (.A0(net284),
    .A1(net148),
    .S(_0584_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(net315),
    .A1(_0596_),
    .S(net99),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _4049_ (.A1(net206),
    .A2(net8),
    .B1(_0568_),
    .B2(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(_0598_),
    .A1(net431),
    .S(_0595_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(\as1802.P[1] ),
    .A1(net238),
    .S(_0584_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _4052_ (.A0(net170),
    .A1(_0599_),
    .S(net99),
    .X(_0600_));
 sky130_fd_sc_hd__o22a_1 _4053_ (.A1(net211),
    .A2(net9),
    .B1(_0569_),
    .B2(net328),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(_0601_),
    .A1(net278),
    .S(_0595_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _4055_ (.A0(net776),
    .A1(net142),
    .S(_0584_),
    .X(_0602_));
 sky130_fd_sc_hd__or2_1 _4056_ (.A(_0513_),
    .B(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__or2_1 _4057_ (.A(net821),
    .B(net99),
    .X(_0604_));
 sky130_fd_sc_hd__a32o_1 _4058_ (.A1(_0568_),
    .A2(_0603_),
    .A3(_0604_),
    .B1(net10),
    .B2(net206),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(_0605_),
    .A1(net819),
    .S(_0595_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(net310),
    .A1(net533),
    .S(_0584_),
    .X(_0606_));
 sky130_fd_sc_hd__or2_1 _4061_ (.A(_0513_),
    .B(net534),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _4062_ (.A(net118),
    .B(_0513_),
    .Y(_0608_));
 sky130_fd_sc_hd__a32o_1 _4063_ (.A1(_0568_),
    .A2(_0607_),
    .A3(_0608_),
    .B1(net11),
    .B2(net206),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(_0609_),
    .A1(net472),
    .S(_0595_),
    .X(_0019_));
 sky130_fd_sc_hd__and3_1 _4065_ (.A(\as1802.instr_latch[7] ),
    .B(net211),
    .C(_0544_),
    .X(_0610_));
 sky130_fd_sc_hd__or4b_1 _4066_ (.A(_3501_),
    .B(_0542_),
    .C(_0581_),
    .D_N(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__or4b_1 _4067_ (.A(_0567_),
    .B(_0577_),
    .C(_0588_),
    .D_N(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__or2_4 _4068_ (.A(_0563_),
    .B(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(net315),
    .A1(net160),
    .S(net99),
    .X(_0614_));
 sky130_fd_sc_hd__o22a_1 _4070_ (.A1(net211),
    .A2(net13),
    .B1(_0569_),
    .B2(net316),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(_0615_),
    .A1(net284),
    .S(_0613_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _4072_ (.A0(net170),
    .A1(net828),
    .S(net99),
    .X(_0616_));
 sky130_fd_sc_hd__a22o_1 _4073_ (.A1(net206),
    .A2(net14),
    .B1(_0568_),
    .B2(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(_0617_),
    .A1(net742),
    .S(_0613_),
    .X(_0021_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(net107),
    .B(net99),
    .Y(_0618_));
 sky130_fd_sc_hd__a32o_1 _4076_ (.A1(_0568_),
    .A2(_0604_),
    .A3(_0618_),
    .B1(net15),
    .B2(net206),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(_0619_),
    .A1(net776),
    .S(_0613_),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _4078_ (.A(net106),
    .B(net99),
    .Y(_0620_));
 sky130_fd_sc_hd__a32o_1 _4079_ (.A1(_0568_),
    .A2(_0608_),
    .A3(_0620_),
    .B1(net16),
    .B2(net206),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _4080_ (.A0(_0621_),
    .A1(net310),
    .S(_0613_),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_8 _4081_ (.A(_0528_),
    .B(_0570_),
    .Y(_0622_));
 sky130_fd_sc_hd__or3_4 _4082_ (.A(net161),
    .B(_0543_),
    .C(_0571_),
    .X(_0623_));
 sky130_fd_sc_hd__and4_4 _4083_ (.A(net161),
    .B(_3496_),
    .C(_0550_),
    .D(_0570_),
    .X(_0624_));
 sky130_fd_sc_hd__nand4_4 _4084_ (.A(net161),
    .B(_3496_),
    .C(_0550_),
    .D(_0570_),
    .Y(_0625_));
 sky130_fd_sc_hd__o21a_4 _4085_ (.A1(_0540_),
    .A2(_0571_),
    .B1(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__and3_2 _4086_ (.A(_0622_),
    .B(_0623_),
    .C(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_2 _4087_ (.A0(net166),
    .A1(net11),
    .S(net83),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_2 _4088_ (.A0(net887),
    .A1(net10),
    .S(net83),
    .X(_0629_));
 sky130_fd_sc_hd__nand2_2 _4089_ (.A(_0628_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__mux2_2 _4090_ (.A0(net170),
    .A1(net9),
    .S(net83),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_4 _4091_ (.A0(\as1802.instr_latch[0] ),
    .A1(net8),
    .S(net83),
    .X(_0632_));
 sky130_fd_sc_hd__nand2_4 _4092_ (.A(_0631_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__and3_2 _4093_ (.A(net212),
    .B(_0623_),
    .C(_0626_),
    .X(_0634_));
 sky130_fd_sc_hd__nand3_4 _4094_ (.A(net212),
    .B(_0623_),
    .C(_0626_),
    .Y(_0635_));
 sky130_fd_sc_hd__or3_4 _4095_ (.A(_0630_),
    .B(_0633_),
    .C(_0634_),
    .X(_0636_));
 sky130_fd_sc_hd__or2_1 _4096_ (.A(_0420_),
    .B(_0428_),
    .X(_0637_));
 sky130_fd_sc_hd__or2_1 _4097_ (.A(_0412_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__or2_1 _4098_ (.A(_0404_),
    .B(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__or2_1 _4099_ (.A(_0396_),
    .B(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__nor2_1 _4100_ (.A(_0388_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_1 _4101_ (.A(_0442_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor2_1 _4102_ (.A(_0451_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _4103_ (.A(_3623_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__o21a_1 _4104_ (.A1(_3623_),
    .A2(_0643_),
    .B1(_0623_),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_4 _4105_ (.A(_3498_),
    .B(_0570_),
    .Y(_0646_));
 sky130_fd_sc_hd__and2_2 _4106_ (.A(_0625_),
    .B(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__nand2_2 _4107_ (.A(_0625_),
    .B(_0646_),
    .Y(_0648_));
 sky130_fd_sc_hd__a2bb2o_1 _4108_ (.A1_N(_3438_),
    .A2_N(_0623_),
    .B1(_0644_),
    .B2(_0645_),
    .X(_0649_));
 sky130_fd_sc_hd__a21o_1 _4109_ (.A1(_3623_),
    .A2(_0452_),
    .B1(_0647_),
    .X(_0650_));
 sky130_fd_sc_hd__o22a_1 _4110_ (.A1(_0648_),
    .A2(_0649_),
    .B1(_0650_),
    .B2(_0453_),
    .X(_0651_));
 sky130_fd_sc_hd__or2_4 _4111_ (.A(net83),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__and3_2 _4112_ (.A(net166),
    .B(_0511_),
    .C(_0570_),
    .X(_0653_));
 sky130_fd_sc_hd__nand3_2 _4113_ (.A(net166),
    .B(_0511_),
    .C(_0570_),
    .Y(_0654_));
 sky130_fd_sc_hd__a32o_1 _4114_ (.A1(_3432_),
    .A2(net171),
    .A3(net96),
    .B1(_3536_),
    .B2(_3537_),
    .X(_0655_));
 sky130_fd_sc_hd__and3_1 _4115_ (.A(net211),
    .B(net104),
    .C(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_2 _4116_ (.A(_0525_),
    .B(_0571_),
    .Y(_0657_));
 sky130_fd_sc_hd__or2_4 _4117_ (.A(_0525_),
    .B(_0571_),
    .X(_0658_));
 sky130_fd_sc_hd__or4_2 _4118_ (.A(_0572_),
    .B(_0653_),
    .C(_0656_),
    .D(net82),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_2 _4119_ (.A(_3498_),
    .B(_0571_),
    .Y(_0660_));
 sky130_fd_sc_hd__and3_2 _4120_ (.A(_3521_),
    .B(_0550_),
    .C(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__nand3_2 _4121_ (.A(_3521_),
    .B(_0550_),
    .C(_0660_),
    .Y(_0662_));
 sky130_fd_sc_hd__or4_4 _4122_ (.A(net173),
    .B(net171),
    .C(_3528_),
    .D(_0509_),
    .X(_0663_));
 sky130_fd_sc_hd__nand2_2 _4123_ (.A(_0662_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__and2b_1 _4124_ (.A_N(_3507_),
    .B(_3520_),
    .X(_0665_));
 sky130_fd_sc_hd__or3b_1 _4125_ (.A(net95),
    .B(_3506_),
    .C_N(_3520_),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _4126_ (.A(net171),
    .B(net211),
    .C(_3494_),
    .X(_0667_));
 sky130_fd_sc_hd__and3_1 _4127_ (.A(_3521_),
    .B(_3552_),
    .C(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _4128_ (.A(_3494_),
    .B(_0570_),
    .C(_0665_),
    .X(_0669_));
 sky130_fd_sc_hd__a21o_1 _4129_ (.A1(_0498_),
    .A2(_0669_),
    .B1(_0668_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _4130_ (.A(\as1802.instr_latch[6] ),
    .B(net171),
    .C(net211),
    .X(_0671_));
 sky130_fd_sc_hd__o2111a_1 _4131_ (.A1(_3492_),
    .A2(_3523_),
    .B1(_0568_),
    .C1(_0665_),
    .D1(_3485_),
    .X(_0672_));
 sky130_fd_sc_hd__nor3_4 _4132_ (.A(_0659_),
    .B(_0664_),
    .C(_0670_),
    .Y(_0673_));
 sky130_fd_sc_hd__and4_4 _4133_ (.A(_3463_),
    .B(\as1802.instr_cycle[1] ),
    .C(_3521_),
    .D(_0660_),
    .X(_0674_));
 sky130_fd_sc_hd__nand4_4 _4134_ (.A(_3463_),
    .B(\as1802.instr_cycle[1] ),
    .C(_3521_),
    .D(_0660_),
    .Y(_0675_));
 sky130_fd_sc_hd__and2_4 _4135_ (.A(_0673_),
    .B(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(_0673_),
    .B(_0675_),
    .Y(_0677_));
 sky130_fd_sc_hd__nor2_2 _4137_ (.A(net172),
    .B(_3525_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _4138_ (.A(_3576_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nor2_2 _4139_ (.A(_0539_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2b_1 _4140_ (.A_N(net169),
    .B(_0515_),
    .Y(_0681_));
 sky130_fd_sc_hd__a32o_1 _4141_ (.A1(_3561_),
    .A2(net99),
    .A3(_0681_),
    .B1(_0542_),
    .B2(net162),
    .X(_0682_));
 sky130_fd_sc_hd__and2_1 _4142_ (.A(_3552_),
    .B(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__o21a_1 _4143_ (.A1(_0680_),
    .A2(_0683_),
    .B1(net211),
    .X(_0684_));
 sky130_fd_sc_hd__o21ai_4 _4144_ (.A1(_0680_),
    .A2(_0683_),
    .B1(net211),
    .Y(_0685_));
 sky130_fd_sc_hd__mux2_1 _4145_ (.A0(\as1802.P[3] ),
    .A1(net16),
    .S(_0676_),
    .X(_0686_));
 sky130_fd_sc_hd__and3_4 _4146_ (.A(net99),
    .B(_0570_),
    .C(net93),
    .X(_0687_));
 sky130_fd_sc_hd__or3_2 _4147_ (.A(_0513_),
    .B(_0571_),
    .C(_0584_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_2 _4148_ (.A0(\as1802.X[3] ),
    .A1(_0686_),
    .S(net80),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(net84),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(\as1802.P[2] ),
    .A1(net15),
    .S(_0676_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_2 _4151_ (.A0(\as1802.X[2] ),
    .A1(_0691_),
    .S(net80),
    .X(_0692_));
 sky130_fd_sc_hd__nand2_1 _4152_ (.A(net84),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__nor2_4 _4153_ (.A(_0690_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(\as1802.P[1] ),
    .A1(net14),
    .S(_0676_),
    .X(_0695_));
 sky130_fd_sc_hd__a21o_1 _4155_ (.A1(\as1802.X[1] ),
    .A2(net81),
    .B1(_0687_),
    .X(_0696_));
 sky130_fd_sc_hd__a21o_2 _4156_ (.A1(net80),
    .A2(_0695_),
    .B1(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__inv_2 _4157_ (.A(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__mux2_1 _4158_ (.A0(\as1802.P[0] ),
    .A1(net13),
    .S(_0676_),
    .X(_0699_));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(\as1802.X[0] ),
    .B(net80),
    .X(_0700_));
 sky130_fd_sc_hd__o211a_2 _4160_ (.A1(net81),
    .A2(_0699_),
    .B1(_0700_),
    .C1(net84),
    .X(_0701_));
 sky130_fd_sc_hd__and2_2 _4161_ (.A(_0697_),
    .B(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__and3_2 _4162_ (.A(net211),
    .B(net80),
    .C(net84),
    .X(_0703_));
 sky130_fd_sc_hd__or4b_4 _4163_ (.A(_0659_),
    .B(_0670_),
    .C(_0674_),
    .D_N(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__and3_4 _4164_ (.A(_0694_),
    .B(_0702_),
    .C(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__or3_2 _4165_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .C(\as1802.regs[2][2] ),
    .X(_0706_));
 sky130_fd_sc_hd__or2_2 _4166_ (.A(\as1802.regs[2][3] ),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__or3_1 _4167_ (.A(\as1802.regs[2][4] ),
    .B(\as1802.regs[2][5] ),
    .C(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__or2_2 _4168_ (.A(\as1802.regs[2][6] ),
    .B(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__nor2_1 _4169_ (.A(\as1802.regs[2][7] ),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__xnor2_1 _4170_ (.A(net840),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__nor2_1 _4171_ (.A(net85),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__mux4_1 _4172_ (.A0(\as1802.regs[8][8] ),
    .A1(\as1802.regs[9][8] ),
    .A2(\as1802.regs[10][8] ),
    .A3(\as1802.regs[11][8] ),
    .S0(net184),
    .S1(net180),
    .X(_0713_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(net113),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__mux4_1 _4174_ (.A0(\as1802.regs[12][8] ),
    .A1(\as1802.regs[13][8] ),
    .A2(\as1802.regs[14][8] ),
    .A3(\as1802.regs[15][8] ),
    .S0(net184),
    .S1(net180),
    .X(_0715_));
 sky130_fd_sc_hd__mux4_1 _4175_ (.A0(\as1802.regs[4][8] ),
    .A1(\as1802.regs[5][8] ),
    .A2(\as1802.regs[6][8] ),
    .A3(\as1802.regs[7][8] ),
    .S0(net184),
    .S1(net180),
    .X(_0716_));
 sky130_fd_sc_hd__mux4_1 _4176_ (.A0(\as1802.regs[0][8] ),
    .A1(\as1802.regs[1][8] ),
    .A2(\as1802.regs[2][8] ),
    .A3(\as1802.regs[3][8] ),
    .S0(net184),
    .S1(net180),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(_0716_),
    .A1(_0717_),
    .S(net113),
    .X(_0718_));
 sky130_fd_sc_hd__a21oi_1 _4178_ (.A1(net176),
    .A2(_0715_),
    .B1(_3470_),
    .Y(_0719_));
 sky130_fd_sc_hd__a2bb2o_2 _4179_ (.A1_N(net175),
    .A2_N(_0718_),
    .B1(_0719_),
    .B2(_0714_),
    .X(_0720_));
 sky130_fd_sc_hd__inv_2 _4180_ (.A(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__mux4_1 _4181_ (.A0(\as1802.regs[12][1] ),
    .A1(\as1802.regs[13][1] ),
    .A2(\as1802.regs[14][1] ),
    .A3(\as1802.regs[15][1] ),
    .S0(net181),
    .S1(net177),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _4182_ (.A(net176),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__mux4_1 _4183_ (.A0(\as1802.regs[8][1] ),
    .A1(\as1802.regs[9][1] ),
    .A2(\as1802.regs[10][1] ),
    .A3(\as1802.regs[11][1] ),
    .S0(net181),
    .S1(net177),
    .X(_0724_));
 sky130_fd_sc_hd__mux4_1 _4184_ (.A0(\as1802.regs[4][1] ),
    .A1(\as1802.regs[5][1] ),
    .A2(\as1802.regs[6][1] ),
    .A3(\as1802.regs[7][1] ),
    .S0(net181),
    .S1(net177),
    .X(_0725_));
 sky130_fd_sc_hd__mux4_1 _4185_ (.A0(\as1802.regs[0][1] ),
    .A1(\as1802.regs[1][1] ),
    .A2(\as1802.regs[2][1] ),
    .A3(\as1802.regs[3][1] ),
    .S0(net181),
    .S1(net177),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _4186_ (.A0(_0725_),
    .A1(_0726_),
    .S(net112),
    .X(_0727_));
 sky130_fd_sc_hd__a21oi_1 _4187_ (.A1(net112),
    .A2(_0724_),
    .B1(_3470_),
    .Y(_0728_));
 sky130_fd_sc_hd__a2bb2o_2 _4188_ (.A1_N(net175),
    .A2_N(_0727_),
    .B1(_0728_),
    .B2(_0723_),
    .X(_0729_));
 sky130_fd_sc_hd__inv_2 _4189_ (.A(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__mux4_1 _4190_ (.A0(\as1802.regs[8][2] ),
    .A1(\as1802.regs[9][2] ),
    .A2(\as1802.regs[10][2] ),
    .A3(\as1802.regs[11][2] ),
    .S0(net182),
    .S1(net178),
    .X(_0731_));
 sky130_fd_sc_hd__mux4_1 _4191_ (.A0(\as1802.regs[12][2] ),
    .A1(\as1802.regs[13][2] ),
    .A2(\as1802.regs[14][2] ),
    .A3(\as1802.regs[15][2] ),
    .S0(net181),
    .S1(net177),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _4192_ (.A(net176),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__mux4_1 _4193_ (.A0(\as1802.regs[4][2] ),
    .A1(\as1802.regs[5][2] ),
    .A2(\as1802.regs[6][2] ),
    .A3(\as1802.regs[7][2] ),
    .S0(net181),
    .S1(net177),
    .X(_0734_));
 sky130_fd_sc_hd__mux4_1 _4194_ (.A0(\as1802.regs[0][2] ),
    .A1(\as1802.regs[1][2] ),
    .A2(\as1802.regs[2][2] ),
    .A3(\as1802.regs[3][2] ),
    .S0(net181),
    .S1(net177),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(_0734_),
    .A1(_0735_),
    .S(net112),
    .X(_0736_));
 sky130_fd_sc_hd__a21oi_1 _4196_ (.A1(net112),
    .A2(_0731_),
    .B1(_3470_),
    .Y(_0737_));
 sky130_fd_sc_hd__a2bb2o_2 _4197_ (.A1_N(net175),
    .A2_N(_0736_),
    .B1(_0737_),
    .B2(_0733_),
    .X(_0738_));
 sky130_fd_sc_hd__inv_2 _4198_ (.A(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_1 _4199_ (.A(_0729_),
    .B(_0738_),
    .Y(_0740_));
 sky130_fd_sc_hd__mux4_1 _4200_ (.A0(\as1802.regs[8][3] ),
    .A1(\as1802.regs[9][3] ),
    .A2(\as1802.regs[10][3] ),
    .A3(\as1802.regs[11][3] ),
    .S0(net182),
    .S1(net178),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_1 _4201_ (.A(net112),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__mux4_1 _4202_ (.A0(\as1802.regs[12][3] ),
    .A1(\as1802.regs[13][3] ),
    .A2(\as1802.regs[14][3] ),
    .A3(\as1802.regs[15][3] ),
    .S0(net181),
    .S1(net177),
    .X(_0743_));
 sky130_fd_sc_hd__mux4_1 _4203_ (.A0(\as1802.regs[4][3] ),
    .A1(\as1802.regs[5][3] ),
    .A2(\as1802.regs[6][3] ),
    .A3(\as1802.regs[7][3] ),
    .S0(net182),
    .S1(net178),
    .X(_0744_));
 sky130_fd_sc_hd__mux4_1 _4204_ (.A0(\as1802.regs[0][3] ),
    .A1(\as1802.regs[1][3] ),
    .A2(\as1802.regs[2][3] ),
    .A3(\as1802.regs[3][3] ),
    .S0(net181),
    .S1(net177),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(_0744_),
    .A1(_0745_),
    .S(net112),
    .X(_0746_));
 sky130_fd_sc_hd__a21oi_1 _4206_ (.A1(net176),
    .A2(_0743_),
    .B1(_3470_),
    .Y(_0747_));
 sky130_fd_sc_hd__a2bb2o_2 _4207_ (.A1_N(net175),
    .A2_N(_0746_),
    .B1(_0747_),
    .B2(_0742_),
    .X(_0748_));
 sky130_fd_sc_hd__inv_2 _4208_ (.A(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__and2_2 _4209_ (.A(_0740_),
    .B(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__mux4_1 _4210_ (.A0(\as1802.regs[8][4] ),
    .A1(\as1802.regs[9][4] ),
    .A2(\as1802.regs[10][4] ),
    .A3(\as1802.regs[11][4] ),
    .S0(net182),
    .S1(net178),
    .X(_0751_));
 sky130_fd_sc_hd__mux4_1 _4211_ (.A0(\as1802.regs[12][4] ),
    .A1(\as1802.regs[13][4] ),
    .A2(\as1802.regs[14][4] ),
    .A3(\as1802.regs[15][4] ),
    .S0(net181),
    .S1(net177),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_1 _4212_ (.A(net176),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__mux4_1 _4213_ (.A0(\as1802.regs[4][4] ),
    .A1(\as1802.regs[5][4] ),
    .A2(\as1802.regs[6][4] ),
    .A3(\as1802.regs[7][4] ),
    .S0(net181),
    .S1(net177),
    .X(_0754_));
 sky130_fd_sc_hd__mux4_1 _4214_ (.A0(\as1802.regs[0][4] ),
    .A1(\as1802.regs[1][4] ),
    .A2(\as1802.regs[2][4] ),
    .A3(\as1802.regs[3][4] ),
    .S0(net181),
    .S1(net177),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(_0754_),
    .A1(_0755_),
    .S(net112),
    .X(_0756_));
 sky130_fd_sc_hd__a21oi_1 _4216_ (.A1(net112),
    .A2(_0751_),
    .B1(_3470_),
    .Y(_0757_));
 sky130_fd_sc_hd__a2bb2o_2 _4217_ (.A1_N(net175),
    .A2_N(_0756_),
    .B1(_0757_),
    .B2(_0753_),
    .X(_0758_));
 sky130_fd_sc_hd__inv_2 _4218_ (.A(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _4219_ (.A(_0750_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__mux4_1 _4220_ (.A0(\as1802.regs[8][5] ),
    .A1(\as1802.regs[9][5] ),
    .A2(\as1802.regs[10][5] ),
    .A3(\as1802.regs[11][5] ),
    .S0(net182),
    .S1(net178),
    .X(_0761_));
 sky130_fd_sc_hd__nand2_1 _4221_ (.A(net112),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__mux4_1 _4222_ (.A0(\as1802.regs[12][5] ),
    .A1(\as1802.regs[13][5] ),
    .A2(\as1802.regs[14][5] ),
    .A3(\as1802.regs[15][5] ),
    .S0(net182),
    .S1(net178),
    .X(_0763_));
 sky130_fd_sc_hd__mux4_1 _4223_ (.A0(\as1802.regs[4][5] ),
    .A1(\as1802.regs[5][5] ),
    .A2(\as1802.regs[6][5] ),
    .A3(\as1802.regs[7][5] ),
    .S0(net182),
    .S1(net178),
    .X(_0764_));
 sky130_fd_sc_hd__mux4_1 _4224_ (.A0(\as1802.regs[0][5] ),
    .A1(\as1802.regs[1][5] ),
    .A2(\as1802.regs[2][5] ),
    .A3(\as1802.regs[3][5] ),
    .S0(net182),
    .S1(net178),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(_0764_),
    .A1(_0765_),
    .S(net112),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_1 _4226_ (.A1(net176),
    .A2(_0763_),
    .B1(_3470_),
    .Y(_0767_));
 sky130_fd_sc_hd__a2bb2o_2 _4227_ (.A1_N(net175),
    .A2_N(_0766_),
    .B1(_0767_),
    .B2(_0762_),
    .X(_0768_));
 sky130_fd_sc_hd__inv_2 _4228_ (.A(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__nor2_1 _4229_ (.A(_0760_),
    .B(_0768_),
    .Y(_0770_));
 sky130_fd_sc_hd__mux4_1 _4230_ (.A0(\as1802.regs[8][6] ),
    .A1(\as1802.regs[9][6] ),
    .A2(\as1802.regs[10][6] ),
    .A3(\as1802.regs[11][6] ),
    .S0(_0008_),
    .S1(_0009_),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_1 _4231_ (.A0(\as1802.regs[12][6] ),
    .A1(\as1802.regs[13][6] ),
    .A2(\as1802.regs[14][6] ),
    .A3(\as1802.regs[15][6] ),
    .S0(net182),
    .S1(net178),
    .X(_0772_));
 sky130_fd_sc_hd__nand2_1 _4232_ (.A(net176),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__mux4_1 _4233_ (.A0(\as1802.regs[4][6] ),
    .A1(\as1802.regs[5][6] ),
    .A2(\as1802.regs[6][6] ),
    .A3(\as1802.regs[7][6] ),
    .S0(net182),
    .S1(net178),
    .X(_0774_));
 sky130_fd_sc_hd__mux4_1 _4234_ (.A0(\as1802.regs[0][6] ),
    .A1(\as1802.regs[1][6] ),
    .A2(\as1802.regs[2][6] ),
    .A3(\as1802.regs[3][6] ),
    .S0(net182),
    .S1(net178),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(_0774_),
    .A1(_0775_),
    .S(net112),
    .X(_0776_));
 sky130_fd_sc_hd__a21oi_1 _4236_ (.A1(net112),
    .A2(_0771_),
    .B1(_3470_),
    .Y(_0777_));
 sky130_fd_sc_hd__a2bb2o_2 _4237_ (.A1_N(net175),
    .A2_N(_0776_),
    .B1(_0777_),
    .B2(_0773_),
    .X(_0778_));
 sky130_fd_sc_hd__inv_2 _4238_ (.A(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _4239_ (.A(_0770_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__mux4_1 _4240_ (.A0(\as1802.regs[8][7] ),
    .A1(\as1802.regs[9][7] ),
    .A2(\as1802.regs[10][7] ),
    .A3(\as1802.regs[11][7] ),
    .S0(net182),
    .S1(net178),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(net112),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__mux4_1 _4242_ (.A0(\as1802.regs[12][7] ),
    .A1(\as1802.regs[13][7] ),
    .A2(\as1802.regs[14][7] ),
    .A3(\as1802.regs[15][7] ),
    .S0(net182),
    .S1(net178),
    .X(_0783_));
 sky130_fd_sc_hd__mux4_1 _4243_ (.A0(\as1802.regs[4][7] ),
    .A1(\as1802.regs[5][7] ),
    .A2(\as1802.regs[6][7] ),
    .A3(\as1802.regs[7][7] ),
    .S0(net182),
    .S1(net178),
    .X(_0784_));
 sky130_fd_sc_hd__mux4_1 _4244_ (.A0(\as1802.regs[0][7] ),
    .A1(\as1802.regs[1][7] ),
    .A2(\as1802.regs[2][7] ),
    .A3(\as1802.regs[3][7] ),
    .S0(net182),
    .S1(net178),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(_0784_),
    .A1(_0785_),
    .S(net113),
    .X(_0786_));
 sky130_fd_sc_hd__a21oi_1 _4246_ (.A1(_0010_),
    .A2(_0783_),
    .B1(_3470_),
    .Y(_0787_));
 sky130_fd_sc_hd__a2bb2o_2 _4247_ (.A1_N(_0011_),
    .A2_N(_0786_),
    .B1(_0787_),
    .B2(_0782_),
    .X(_0788_));
 sky130_fd_sc_hd__inv_2 _4248_ (.A(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(_0780_),
    .B(_0788_),
    .X(_0790_));
 sky130_fd_sc_hd__or2_1 _4250_ (.A(_0720_),
    .B(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__mux4_1 _4251_ (.A0(\as1802.regs[8][0] ),
    .A1(\as1802.regs[9][0] ),
    .A2(\as1802.regs[10][0] ),
    .A3(\as1802.regs[11][0] ),
    .S0(net181),
    .S1(net177),
    .X(_0792_));
 sky130_fd_sc_hd__mux4_1 _4252_ (.A0(\as1802.regs[12][0] ),
    .A1(\as1802.regs[13][0] ),
    .A2(\as1802.regs[14][0] ),
    .A3(\as1802.regs[15][0] ),
    .S0(net181),
    .S1(net177),
    .X(_0793_));
 sky130_fd_sc_hd__or2_1 _4253_ (.A(net112),
    .B(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__mux4_1 _4254_ (.A0(\as1802.regs[4][0] ),
    .A1(\as1802.regs[5][0] ),
    .A2(\as1802.regs[6][0] ),
    .A3(\as1802.regs[7][0] ),
    .S0(net181),
    .S1(net177),
    .X(_0795_));
 sky130_fd_sc_hd__mux4_1 _4255_ (.A0(\as1802.regs[0][0] ),
    .A1(\as1802.regs[1][0] ),
    .A2(\as1802.regs[2][0] ),
    .A3(\as1802.regs[3][0] ),
    .S0(net181),
    .S1(net177),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(_0795_),
    .A1(_0796_),
    .S(net112),
    .X(_0797_));
 sky130_fd_sc_hd__o211a_1 _4257_ (.A1(net176),
    .A2(_0792_),
    .B1(_0794_),
    .C1(net175),
    .X(_0798_));
 sky130_fd_sc_hd__a21oi_4 _4258_ (.A1(_3470_),
    .A2(_0797_),
    .B1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__inv_2 _4259_ (.A(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__or2_1 _4260_ (.A(_0791_),
    .B(_0799_),
    .X(_0801_));
 sky130_fd_sc_hd__nor2_1 _4261_ (.A(_0790_),
    .B(_0799_),
    .Y(_0802_));
 sky130_fd_sc_hd__o21a_1 _4262_ (.A1(_0721_),
    .A2(_0802_),
    .B1(_0801_),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_1 _4263_ (.A(net165),
    .B(_0573_),
    .Y(_0804_));
 sky130_fd_sc_hd__mux2_2 _4264_ (.A0(_0668_),
    .A1(_0669_),
    .S(_0498_),
    .X(_0805_));
 sky130_fd_sc_hd__inv_2 _4265_ (.A(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__nor2_1 _4266_ (.A(_0804_),
    .B(_0805_),
    .Y(_0807_));
 sky130_fd_sc_hd__and4b_1 _4267_ (.A_N(_0498_),
    .B(_0671_),
    .C(_3521_),
    .D(_3552_),
    .X(_0808_));
 sky130_fd_sc_hd__a31o_2 _4268_ (.A1(_0498_),
    .A2(_0541_),
    .A3(_0672_),
    .B1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__or2_2 _4269_ (.A(_0804_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__or2_1 _4270_ (.A(net165),
    .B(_0720_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _4271_ (.A(_0720_),
    .B(_0790_),
    .Y(_0812_));
 sky130_fd_sc_hd__nand3_1 _4272_ (.A(_0791_),
    .B(_0809_),
    .C(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__o2bb2a_1 _4273_ (.A1_N(_0803_),
    .A2_N(_0807_),
    .B1(_0811_),
    .B2(_0573_),
    .X(_0814_));
 sky130_fd_sc_hd__a21oi_1 _4274_ (.A1(_0813_),
    .A2(_0814_),
    .B1(_0674_),
    .Y(_0815_));
 sky130_fd_sc_hd__a211o_1 _4275_ (.A1(net160),
    .A2(_0674_),
    .B1(_0815_),
    .C1(net82),
    .X(_0816_));
 sky130_fd_sc_hd__a21bo_1 _4276_ (.A1(net165),
    .A2(_0803_),
    .B1_N(_0811_),
    .X(_0817_));
 sky130_fd_sc_hd__o211a_1 _4277_ (.A1(_0658_),
    .A2(_0817_),
    .B1(_0816_),
    .C1(net78),
    .X(_0818_));
 sky130_fd_sc_hd__a211o_1 _4278_ (.A1(net29),
    .A2(_0676_),
    .B1(_0684_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__and3_4 _4279_ (.A(net162),
    .B(_0542_),
    .C(_0570_),
    .X(_0820_));
 sky130_fd_sc_hd__or3_4 _4280_ (.A(net119),
    .B(_0543_),
    .C(_0571_),
    .X(_0821_));
 sky130_fd_sc_hd__mux4_1 _4281_ (.A0(\as1802.regs[8][8] ),
    .A1(\as1802.regs[9][8] ),
    .A2(\as1802.regs[10][8] ),
    .A3(\as1802.regs[11][8] ),
    .S0(net204),
    .S1(net200),
    .X(_0822_));
 sky130_fd_sc_hd__mux4_1 _4282_ (.A0(\as1802.regs[12][8] ),
    .A1(\as1802.regs[13][8] ),
    .A2(\as1802.regs[14][8] ),
    .A3(\as1802.regs[15][8] ),
    .S0(net204),
    .S1(net200),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(_0822_),
    .A1(_0823_),
    .S(net196),
    .X(_0824_));
 sky130_fd_sc_hd__mux4_1 _4284_ (.A0(\as1802.regs[4][8] ),
    .A1(\as1802.regs[5][8] ),
    .A2(\as1802.regs[6][8] ),
    .A3(\as1802.regs[7][8] ),
    .S0(net205),
    .S1(net201),
    .X(_0825_));
 sky130_fd_sc_hd__mux4_1 _4285_ (.A0(\as1802.regs[0][8] ),
    .A1(\as1802.regs[1][8] ),
    .A2(\as1802.regs[2][8] ),
    .A3(\as1802.regs[3][8] ),
    .S0(net205),
    .S1(net201),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(_0826_),
    .A1(_0825_),
    .S(net196),
    .X(_0827_));
 sky130_fd_sc_hd__and2b_1 _4287_ (.A_N(net194),
    .B(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__a21oi_4 _4288_ (.A1(net194),
    .A2(_0824_),
    .B1(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__or4_2 _4289_ (.A(_3512_),
    .B(_3562_),
    .C(_0513_),
    .D(_0571_),
    .X(_0830_));
 sky130_fd_sc_hd__or4_2 _4290_ (.A(_3512_),
    .B(_3562_),
    .C(_0513_),
    .D(_0571_),
    .X(_0831_));
 sky130_fd_sc_hd__xor2_1 _4291_ (.A(_0829_),
    .B(net90),
    .X(_0832_));
 sky130_fd_sc_hd__mux4_1 _4292_ (.A0(\as1802.regs[8][5] ),
    .A1(\as1802.regs[9][5] ),
    .A2(\as1802.regs[10][5] ),
    .A3(\as1802.regs[11][5] ),
    .S0(net202),
    .S1(net198),
    .X(_0833_));
 sky130_fd_sc_hd__mux4_1 _4293_ (.A0(\as1802.regs[12][5] ),
    .A1(\as1802.regs[13][5] ),
    .A2(\as1802.regs[14][5] ),
    .A3(\as1802.regs[15][5] ),
    .S0(net202),
    .S1(net198),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(_0833_),
    .A1(_0834_),
    .S(net197),
    .X(_0835_));
 sky130_fd_sc_hd__mux4_1 _4295_ (.A0(\as1802.regs[4][5] ),
    .A1(\as1802.regs[5][5] ),
    .A2(\as1802.regs[6][5] ),
    .A3(\as1802.regs[7][5] ),
    .S0(net202),
    .S1(net198),
    .X(_0836_));
 sky130_fd_sc_hd__mux4_1 _4296_ (.A0(\as1802.regs[0][5] ),
    .A1(\as1802.regs[1][5] ),
    .A2(\as1802.regs[2][5] ),
    .A3(\as1802.regs[3][5] ),
    .S0(net203),
    .S1(net199),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(_0837_),
    .A1(_0836_),
    .S(net197),
    .X(_0838_));
 sky130_fd_sc_hd__and2b_1 _4298_ (.A_N(net195),
    .B(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__a21oi_4 _4299_ (.A1(net195),
    .A2(_0835_),
    .B1(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__xnor2_1 _4300_ (.A(net89),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__mux4_1 _4301_ (.A0(\as1802.regs[8][4] ),
    .A1(\as1802.regs[9][4] ),
    .A2(\as1802.regs[10][4] ),
    .A3(\as1802.regs[11][4] ),
    .S0(net202),
    .S1(net198),
    .X(_0842_));
 sky130_fd_sc_hd__mux4_1 _4302_ (.A0(\as1802.regs[12][4] ),
    .A1(\as1802.regs[13][4] ),
    .A2(\as1802.regs[14][4] ),
    .A3(\as1802.regs[15][4] ),
    .S0(net202),
    .S1(net198),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _4303_ (.A0(_0842_),
    .A1(_0843_),
    .S(net197),
    .X(_0844_));
 sky130_fd_sc_hd__nand2b_1 _4304_ (.A_N(_0844_),
    .B(net195),
    .Y(_0845_));
 sky130_fd_sc_hd__mux4_1 _4305_ (.A0(\as1802.regs[4][4] ),
    .A1(\as1802.regs[5][4] ),
    .A2(\as1802.regs[6][4] ),
    .A3(\as1802.regs[7][4] ),
    .S0(net203),
    .S1(net199),
    .X(_0846_));
 sky130_fd_sc_hd__mux4_1 _4306_ (.A0(\as1802.regs[0][4] ),
    .A1(\as1802.regs[1][4] ),
    .A2(\as1802.regs[2][4] ),
    .A3(\as1802.regs[3][4] ),
    .S0(net203),
    .S1(net199),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(_0847_),
    .A1(_0846_),
    .S(net197),
    .X(_0848_));
 sky130_fd_sc_hd__o21ai_4 _4308_ (.A1(net195),
    .A2(_0848_),
    .B1(_0845_),
    .Y(_0849_));
 sky130_fd_sc_hd__and2_1 _4309_ (.A(net89),
    .B(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__nor2_1 _4310_ (.A(net89),
    .B(_0849_),
    .Y(_0851_));
 sky130_fd_sc_hd__or2_1 _4311_ (.A(_0850_),
    .B(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__mux4_1 _4312_ (.A0(\as1802.regs[8][3] ),
    .A1(\as1802.regs[9][3] ),
    .A2(\as1802.regs[10][3] ),
    .A3(\as1802.regs[11][3] ),
    .S0(net202),
    .S1(net198),
    .X(_0853_));
 sky130_fd_sc_hd__mux4_1 _4313_ (.A0(\as1802.regs[12][3] ),
    .A1(\as1802.regs[13][3] ),
    .A2(\as1802.regs[14][3] ),
    .A3(\as1802.regs[15][3] ),
    .S0(net202),
    .S1(net198),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(_0853_),
    .A1(_0854_),
    .S(net197),
    .X(_0855_));
 sky130_fd_sc_hd__mux4_1 _4315_ (.A0(\as1802.regs[4][3] ),
    .A1(\as1802.regs[5][3] ),
    .A2(\as1802.regs[6][3] ),
    .A3(\as1802.regs[7][3] ),
    .S0(net202),
    .S1(net198),
    .X(_0856_));
 sky130_fd_sc_hd__mux4_1 _4316_ (.A0(\as1802.regs[0][3] ),
    .A1(\as1802.regs[1][3] ),
    .A2(\as1802.regs[2][3] ),
    .A3(\as1802.regs[3][3] ),
    .S0(net203),
    .S1(net199),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(_0857_),
    .A1(_0856_),
    .S(net197),
    .X(_0858_));
 sky130_fd_sc_hd__and2b_1 _4318_ (.A_N(net195),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__a21oi_2 _4319_ (.A1(net195),
    .A2(_0855_),
    .B1(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__or2_1 _4320_ (.A(_0830_),
    .B(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__and2_1 _4321_ (.A(net89),
    .B(_0860_),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(net89),
    .B(_0860_),
    .Y(_0863_));
 sky130_fd_sc_hd__mux4_1 _4323_ (.A0(\as1802.regs[8][2] ),
    .A1(\as1802.regs[9][2] ),
    .A2(\as1802.regs[10][2] ),
    .A3(\as1802.regs[11][2] ),
    .S0(net202),
    .S1(net198),
    .X(_0864_));
 sky130_fd_sc_hd__mux4_1 _4324_ (.A0(\as1802.regs[12][2] ),
    .A1(\as1802.regs[13][2] ),
    .A2(\as1802.regs[14][2] ),
    .A3(\as1802.regs[15][2] ),
    .S0(net202),
    .S1(net198),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(_0864_),
    .A1(_0865_),
    .S(net197),
    .X(_0866_));
 sky130_fd_sc_hd__nand2b_1 _4326_ (.A_N(_0866_),
    .B(net195),
    .Y(_0867_));
 sky130_fd_sc_hd__mux4_1 _4327_ (.A0(\as1802.regs[4][2] ),
    .A1(\as1802.regs[5][2] ),
    .A2(\as1802.regs[6][2] ),
    .A3(\as1802.regs[7][2] ),
    .S0(net203),
    .S1(net199),
    .X(_0868_));
 sky130_fd_sc_hd__mux4_1 _4328_ (.A0(\as1802.regs[0][2] ),
    .A1(\as1802.regs[1][2] ),
    .A2(\as1802.regs[2][2] ),
    .A3(\as1802.regs[3][2] ),
    .S0(net203),
    .S1(net199),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(_0869_),
    .A1(_0868_),
    .S(net197),
    .X(_0870_));
 sky130_fd_sc_hd__o21ai_2 _4330_ (.A1(net195),
    .A2(_0870_),
    .B1(_0867_),
    .Y(_0871_));
 sky130_fd_sc_hd__xor2_1 _4331_ (.A(net89),
    .B(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__mux4_1 _4332_ (.A0(\as1802.regs[8][1] ),
    .A1(\as1802.regs[9][1] ),
    .A2(\as1802.regs[10][1] ),
    .A3(\as1802.regs[11][1] ),
    .S0(net202),
    .S1(net198),
    .X(_0873_));
 sky130_fd_sc_hd__mux4_1 _4333_ (.A0(\as1802.regs[12][1] ),
    .A1(\as1802.regs[13][1] ),
    .A2(\as1802.regs[14][1] ),
    .A3(\as1802.regs[15][1] ),
    .S0(net202),
    .S1(net198),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(_0873_),
    .A1(_0874_),
    .S(net197),
    .X(_0875_));
 sky130_fd_sc_hd__nand2b_1 _4335_ (.A_N(_0875_),
    .B(net195),
    .Y(_0876_));
 sky130_fd_sc_hd__mux4_1 _4336_ (.A0(\as1802.regs[4][1] ),
    .A1(\as1802.regs[5][1] ),
    .A2(\as1802.regs[6][1] ),
    .A3(\as1802.regs[7][1] ),
    .S0(net203),
    .S1(net199),
    .X(_0877_));
 sky130_fd_sc_hd__mux4_1 _4337_ (.A0(\as1802.regs[0][1] ),
    .A1(\as1802.regs[1][1] ),
    .A2(\as1802.regs[2][1] ),
    .A3(\as1802.regs[3][1] ),
    .S0(net203),
    .S1(net199),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(_0878_),
    .A1(_0877_),
    .S(net197),
    .X(_0879_));
 sky130_fd_sc_hd__o21ai_2 _4339_ (.A1(net195),
    .A2(_0879_),
    .B1(_0876_),
    .Y(_0880_));
 sky130_fd_sc_hd__xnor2_1 _4340_ (.A(net89),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__mux4_1 _4341_ (.A0(\as1802.regs[8][0] ),
    .A1(\as1802.regs[9][0] ),
    .A2(\as1802.regs[10][0] ),
    .A3(\as1802.regs[11][0] ),
    .S0(net202),
    .S1(net198),
    .X(_0882_));
 sky130_fd_sc_hd__mux4_1 _4342_ (.A0(\as1802.regs[12][0] ),
    .A1(\as1802.regs[13][0] ),
    .A2(\as1802.regs[14][0] ),
    .A3(\as1802.regs[15][0] ),
    .S0(net202),
    .S1(net198),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(_0882_),
    .A1(_0883_),
    .S(net197),
    .X(_0884_));
 sky130_fd_sc_hd__nand2b_1 _4344_ (.A_N(_0884_),
    .B(net195),
    .Y(_0885_));
 sky130_fd_sc_hd__mux4_1 _4345_ (.A0(\as1802.regs[4][0] ),
    .A1(\as1802.regs[5][0] ),
    .A2(\as1802.regs[6][0] ),
    .A3(\as1802.regs[7][0] ),
    .S0(net203),
    .S1(net199),
    .X(_0886_));
 sky130_fd_sc_hd__mux4_1 _4346_ (.A0(\as1802.regs[0][0] ),
    .A1(\as1802.regs[1][0] ),
    .A2(\as1802.regs[2][0] ),
    .A3(\as1802.regs[3][0] ),
    .S0(net203),
    .S1(net199),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(_0887_),
    .A1(_0886_),
    .S(net197),
    .X(_0888_));
 sky130_fd_sc_hd__o21ai_2 _4348_ (.A1(net195),
    .A2(_0888_),
    .B1(_0885_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _4349_ (.A(_0881_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__o21bai_1 _4350_ (.A1(net89),
    .A2(_0880_),
    .B1_N(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__and2_1 _4351_ (.A(_0872_),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__o21ba_1 _4352_ (.A1(net89),
    .A2(_0871_),
    .B1_N(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__nand2_1 _4353_ (.A(_0861_),
    .B(_0863_),
    .Y(_0894_));
 sky130_fd_sc_hd__o21a_1 _4354_ (.A1(_0862_),
    .A2(_0893_),
    .B1(_0861_),
    .X(_0895_));
 sky130_fd_sc_hd__or2_1 _4355_ (.A(_0852_),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__or2_1 _4356_ (.A(_0841_),
    .B(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__mux4_1 _4357_ (.A0(\as1802.regs[8][6] ),
    .A1(\as1802.regs[9][6] ),
    .A2(\as1802.regs[10][6] ),
    .A3(\as1802.regs[11][6] ),
    .S0(net202),
    .S1(net198),
    .X(_0898_));
 sky130_fd_sc_hd__mux4_1 _4358_ (.A0(\as1802.regs[12][6] ),
    .A1(\as1802.regs[13][6] ),
    .A2(\as1802.regs[14][6] ),
    .A3(\as1802.regs[15][6] ),
    .S0(net203),
    .S1(net199),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(_0898_),
    .A1(_0899_),
    .S(net197),
    .X(_0900_));
 sky130_fd_sc_hd__nand2b_1 _4360_ (.A_N(_0900_),
    .B(net195),
    .Y(_0901_));
 sky130_fd_sc_hd__mux4_1 _4361_ (.A0(\as1802.regs[4][6] ),
    .A1(\as1802.regs[5][6] ),
    .A2(\as1802.regs[6][6] ),
    .A3(\as1802.regs[7][6] ),
    .S0(net203),
    .S1(net199),
    .X(_0902_));
 sky130_fd_sc_hd__mux4_1 _4362_ (.A0(\as1802.regs[0][6] ),
    .A1(\as1802.regs[1][6] ),
    .A2(\as1802.regs[2][6] ),
    .A3(\as1802.regs[3][6] ),
    .S0(net203),
    .S1(net199),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _4363_ (.A0(_0903_),
    .A1(_0902_),
    .S(net197),
    .X(_0904_));
 sky130_fd_sc_hd__o21ai_2 _4364_ (.A1(net195),
    .A2(_0904_),
    .B1(_0901_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(net89),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__or2_1 _4366_ (.A(net89),
    .B(_0905_),
    .X(_0907_));
 sky130_fd_sc_hd__nand2_1 _4367_ (.A(_0906_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__mux4_1 _4368_ (.A0(\as1802.regs[8][7] ),
    .A1(\as1802.regs[9][7] ),
    .A2(\as1802.regs[10][7] ),
    .A3(\as1802.regs[11][7] ),
    .S0(net203),
    .S1(net199),
    .X(_0909_));
 sky130_fd_sc_hd__mux4_1 _4369_ (.A0(\as1802.regs[12][7] ),
    .A1(\as1802.regs[13][7] ),
    .A2(\as1802.regs[14][7] ),
    .A3(\as1802.regs[15][7] ),
    .S0(net203),
    .S1(net199),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(_0909_),
    .A1(_0910_),
    .S(_0006_),
    .X(_0911_));
 sky130_fd_sc_hd__mux4_1 _4371_ (.A0(\as1802.regs[4][7] ),
    .A1(\as1802.regs[5][7] ),
    .A2(\as1802.regs[6][7] ),
    .A3(\as1802.regs[7][7] ),
    .S0(net202),
    .S1(net198),
    .X(_0912_));
 sky130_fd_sc_hd__mux4_1 _4372_ (.A0(\as1802.regs[0][7] ),
    .A1(\as1802.regs[1][7] ),
    .A2(\as1802.regs[2][7] ),
    .A3(\as1802.regs[3][7] ),
    .S0(net204),
    .S1(net200),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(_0913_),
    .A1(_0912_),
    .S(net196),
    .X(_0914_));
 sky130_fd_sc_hd__and2b_1 _4374_ (.A_N(net194),
    .B(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a21oi_4 _4375_ (.A1(net194),
    .A2(_0911_),
    .B1(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__xnor2_2 _4376_ (.A(net90),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a41o_1 _4377_ (.A1(_0840_),
    .A2(_0849_),
    .A3(_0905_),
    .A4(_0916_),
    .B1(_0830_),
    .X(_0918_));
 sky130_fd_sc_hd__o31ai_2 _4378_ (.A1(_0897_),
    .A2(_0908_),
    .A3(_0917_),
    .B1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__a21o_1 _4379_ (.A1(_0840_),
    .A2(_0849_),
    .B1(net89),
    .X(_0920_));
 sky130_fd_sc_hd__a31o_1 _4380_ (.A1(_0840_),
    .A2(_0849_),
    .A3(_0916_),
    .B1(net89),
    .X(_0921_));
 sky130_fd_sc_hd__o311a_1 _4381_ (.A1(_0897_),
    .A2(_0908_),
    .A3(_0917_),
    .B1(_0921_),
    .C1(_0907_),
    .X(_0922_));
 sky130_fd_sc_hd__o21a_1 _4382_ (.A1(_0832_),
    .A2(_0919_),
    .B1(_0821_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _4383_ (.A(_0832_),
    .B(_0919_),
    .Y(_0924_));
 sky130_fd_sc_hd__a221o_1 _4384_ (.A1(_3623_),
    .A2(_0820_),
    .B1(_0923_),
    .B2(_0924_),
    .C1(net80),
    .X(_0925_));
 sky130_fd_sc_hd__a31o_4 _4385_ (.A1(net85),
    .A2(_0819_),
    .A3(_0925_),
    .B1(_0712_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _4386_ (.A0(net639),
    .A1(_0926_),
    .S(_0705_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _4387_ (.A0(_0652_),
    .A1(net640),
    .S(_0636_),
    .X(_0028_));
 sky130_fd_sc_hd__or2_1 _4388_ (.A(_3616_),
    .B(_0644_),
    .X(_0928_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_3616_),
    .B(_0644_),
    .Y(_0929_));
 sky130_fd_sc_hd__and3_1 _4390_ (.A(_0623_),
    .B(_0928_),
    .C(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__nor2_1 _4391_ (.A(_3437_),
    .B(_0623_),
    .Y(_0931_));
 sky130_fd_sc_hd__o21ai_1 _4392_ (.A1(_3616_),
    .A2(_0453_),
    .B1(_0648_),
    .Y(_0932_));
 sky130_fd_sc_hd__o32a_1 _4393_ (.A1(_0648_),
    .A2(_0930_),
    .A3(_0931_),
    .B1(_0932_),
    .B2(_0454_),
    .X(_0933_));
 sky130_fd_sc_hd__or2_4 _4394_ (.A(net83),
    .B(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__mux4_1 _4395_ (.A0(\as1802.regs[8][9] ),
    .A1(\as1802.regs[9][9] ),
    .A2(\as1802.regs[10][9] ),
    .A3(\as1802.regs[11][9] ),
    .S0(net184),
    .S1(net180),
    .X(_0935_));
 sky130_fd_sc_hd__mux4_1 _4396_ (.A0(\as1802.regs[12][9] ),
    .A1(\as1802.regs[13][9] ),
    .A2(\as1802.regs[14][9] ),
    .A3(\as1802.regs[15][9] ),
    .S0(net184),
    .S1(net180),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _4397_ (.A0(_0935_),
    .A1(_0936_),
    .S(net176),
    .X(_0937_));
 sky130_fd_sc_hd__and2_1 _4398_ (.A(net175),
    .B(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__mux4_1 _4399_ (.A0(\as1802.regs[4][9] ),
    .A1(\as1802.regs[5][9] ),
    .A2(\as1802.regs[6][9] ),
    .A3(\as1802.regs[7][9] ),
    .S0(net184),
    .S1(net180),
    .X(_0939_));
 sky130_fd_sc_hd__mux4_1 _4400_ (.A0(\as1802.regs[0][9] ),
    .A1(\as1802.regs[1][9] ),
    .A2(\as1802.regs[2][9] ),
    .A3(\as1802.regs[3][9] ),
    .S0(net184),
    .S1(net180),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_1 _4401_ (.A0(_0939_),
    .A1(_0940_),
    .S(net112),
    .X(_0941_));
 sky130_fd_sc_hd__a21oi_4 _4402_ (.A1(_3470_),
    .A2(_0941_),
    .B1(_0938_),
    .Y(_0942_));
 sky130_fd_sc_hd__inv_2 _4403_ (.A(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(_0791_),
    .B(_0942_),
    .X(_0944_));
 sky130_fd_sc_hd__or2_1 _4405_ (.A(_0799_),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__a21bo_1 _4406_ (.A1(_0801_),
    .A2(_0942_),
    .B1_N(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__nand2_1 _4407_ (.A(_0791_),
    .B(_0942_),
    .Y(_0947_));
 sky130_fd_sc_hd__and3_1 _4408_ (.A(_0805_),
    .B(_0944_),
    .C(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__a211o_1 _4409_ (.A1(_0804_),
    .A2(_0943_),
    .B1(_0948_),
    .C1(_0674_),
    .X(_0949_));
 sky130_fd_sc_hd__o21ba_1 _4410_ (.A1(_0810_),
    .A2(_0946_),
    .B1_N(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__a211o_1 _4411_ (.A1(net108),
    .A2(_0674_),
    .B1(_0950_),
    .C1(net82),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(_0942_),
    .A1(_0946_),
    .S(net165),
    .X(_0952_));
 sky130_fd_sc_hd__or2_1 _4413_ (.A(_0658_),
    .B(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__o21ai_1 _4414_ (.A1(net30),
    .A2(net78),
    .B1(net80),
    .Y(_0954_));
 sky130_fd_sc_hd__a31o_1 _4415_ (.A1(net78),
    .A2(_0951_),
    .A3(_0953_),
    .B1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__mux4_1 _4416_ (.A0(\as1802.regs[8][9] ),
    .A1(\as1802.regs[9][9] ),
    .A2(\as1802.regs[10][9] ),
    .A3(\as1802.regs[11][9] ),
    .S0(net204),
    .S1(net200),
    .X(_0956_));
 sky130_fd_sc_hd__mux4_1 _4417_ (.A0(\as1802.regs[12][9] ),
    .A1(\as1802.regs[13][9] ),
    .A2(\as1802.regs[14][9] ),
    .A3(\as1802.regs[15][9] ),
    .S0(net204),
    .S1(net200),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _4418_ (.A0(_0956_),
    .A1(_0957_),
    .S(net196),
    .X(_0958_));
 sky130_fd_sc_hd__mux4_1 _4419_ (.A0(\as1802.regs[4][9] ),
    .A1(\as1802.regs[5][9] ),
    .A2(\as1802.regs[6][9] ),
    .A3(\as1802.regs[7][9] ),
    .S0(net204),
    .S1(net200),
    .X(_0959_));
 sky130_fd_sc_hd__mux4_1 _4420_ (.A0(\as1802.regs[0][9] ),
    .A1(\as1802.regs[1][9] ),
    .A2(\as1802.regs[2][9] ),
    .A3(\as1802.regs[3][9] ),
    .S0(net205),
    .S1(net201),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(_0960_),
    .A1(_0959_),
    .S(net197),
    .X(_0961_));
 sky130_fd_sc_hd__and2b_1 _4422_ (.A_N(net194),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__a21oi_2 _4423_ (.A1(net194),
    .A2(_0958_),
    .B1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__and2_1 _4424_ (.A(net90),
    .B(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__nor2_1 _4425_ (.A(net90),
    .B(_0963_),
    .Y(_0965_));
 sky130_fd_sc_hd__nor2_1 _4426_ (.A(_0964_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__o21a_1 _4427_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0924_),
    .X(_0967_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_0966_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__o21a_1 _4429_ (.A1(_0966_),
    .A2(_0967_),
    .B1(_0821_),
    .X(_0969_));
 sky130_fd_sc_hd__a221o_1 _4430_ (.A1(_3616_),
    .A2(_0820_),
    .B1(_0968_),
    .B2(_0969_),
    .C1(net80),
    .X(_0970_));
 sky130_fd_sc_hd__and3_1 _4431_ (.A(net84),
    .B(_0955_),
    .C(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__or4_4 _4432_ (.A(\as1802.regs[2][7] ),
    .B(\as1802.regs[2][8] ),
    .C(\as1802.regs[2][9] ),
    .D(_0709_),
    .X(_0972_));
 sky130_fd_sc_hd__o31ai_2 _4433_ (.A1(\as1802.regs[2][7] ),
    .A2(\as1802.regs[2][8] ),
    .A3(_0709_),
    .B1(\as1802.regs[2][9] ),
    .Y(_0973_));
 sky130_fd_sc_hd__a31oi_4 _4434_ (.A1(_0687_),
    .A2(_0972_),
    .A3(_0973_),
    .B1(_0971_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(net752),
    .A1(_0974_),
    .S(_0705_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _4436_ (.A0(_0934_),
    .A1(_0975_),
    .S(_0636_),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _4437_ (.A(_0462_),
    .B(_0928_),
    .Y(_0976_));
 sky130_fd_sc_hd__and2_1 _4438_ (.A(_0462_),
    .B(_0928_),
    .X(_0977_));
 sky130_fd_sc_hd__nor2_1 _4439_ (.A(_0976_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__nand2_2 _4440_ (.A(_0623_),
    .B(_0646_),
    .Y(_0979_));
 sky130_fd_sc_hd__o22a_1 _4441_ (.A1(net132),
    .A2(_0623_),
    .B1(_0978_),
    .B2(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__o2bb2a_1 _4442_ (.A1_N(_0488_),
    .A2_N(_0648_),
    .B1(_0980_),
    .B2(_0624_),
    .X(_0981_));
 sky130_fd_sc_hd__or2_4 _4443_ (.A(net83),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__xnor2_1 _4444_ (.A(net874),
    .B(_0972_),
    .Y(_0983_));
 sky130_fd_sc_hd__mux4_1 _4445_ (.A0(\as1802.regs[8][10] ),
    .A1(\as1802.regs[9][10] ),
    .A2(\as1802.regs[10][10] ),
    .A3(\as1802.regs[11][10] ),
    .S0(net184),
    .S1(net180),
    .X(_0984_));
 sky130_fd_sc_hd__mux4_1 _4446_ (.A0(\as1802.regs[12][10] ),
    .A1(\as1802.regs[13][10] ),
    .A2(\as1802.regs[14][10] ),
    .A3(\as1802.regs[15][10] ),
    .S0(net184),
    .S1(net180),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _4447_ (.A0(_0984_),
    .A1(_0985_),
    .S(net176),
    .X(_0986_));
 sky130_fd_sc_hd__and2_1 _4448_ (.A(net175),
    .B(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__mux4_1 _4449_ (.A0(\as1802.regs[4][10] ),
    .A1(\as1802.regs[5][10] ),
    .A2(\as1802.regs[6][10] ),
    .A3(\as1802.regs[7][10] ),
    .S0(net184),
    .S1(net180),
    .X(_0988_));
 sky130_fd_sc_hd__mux4_1 _4450_ (.A0(\as1802.regs[0][10] ),
    .A1(\as1802.regs[1][10] ),
    .A2(\as1802.regs[2][10] ),
    .A3(\as1802.regs[3][10] ),
    .S0(net184),
    .S1(net180),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(_0988_),
    .A1(_0989_),
    .S(net113),
    .X(_0990_));
 sky130_fd_sc_hd__a21oi_4 _4452_ (.A1(_3470_),
    .A2(_0990_),
    .B1(_0987_),
    .Y(_0991_));
 sky130_fd_sc_hd__inv_2 _4453_ (.A(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__or2_1 _4454_ (.A(_0944_),
    .B(_0991_),
    .X(_0993_));
 sky130_fd_sc_hd__o2bb2a_1 _4455_ (.A1_N(_0945_),
    .A2_N(_0991_),
    .B1(_0993_),
    .B2(_0799_),
    .X(_0994_));
 sky130_fd_sc_hd__o21ai_1 _4456_ (.A1(_0806_),
    .A2(_0944_),
    .B1(_0991_),
    .Y(_0995_));
 sky130_fd_sc_hd__o21a_1 _4457_ (.A1(_0806_),
    .A2(_0993_),
    .B1(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(_0994_),
    .A1(_0996_),
    .S(_0810_),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(net154),
    .A1(_0997_),
    .S(_0675_),
    .X(_0998_));
 sky130_fd_sc_hd__nor2_1 _4460_ (.A(net165),
    .B(_0991_),
    .Y(_0999_));
 sky130_fd_sc_hd__a211o_1 _4461_ (.A1(net165),
    .A2(_0994_),
    .B1(_0999_),
    .C1(_0658_),
    .X(_1000_));
 sky130_fd_sc_hd__o211a_1 _4462_ (.A1(_0657_),
    .A2(_0998_),
    .B1(_1000_),
    .C1(_0654_),
    .X(_1001_));
 sky130_fd_sc_hd__a21o_1 _4463_ (.A1(_0653_),
    .A2(_0994_),
    .B1(_0676_),
    .X(_1002_));
 sky130_fd_sc_hd__o22a_1 _4464_ (.A1(net2),
    .A2(net78),
    .B1(_1001_),
    .B2(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__mux4_1 _4465_ (.A0(\as1802.regs[8][10] ),
    .A1(\as1802.regs[9][10] ),
    .A2(\as1802.regs[10][10] ),
    .A3(\as1802.regs[11][10] ),
    .S0(net204),
    .S1(net200),
    .X(_1004_));
 sky130_fd_sc_hd__mux4_1 _4466_ (.A0(\as1802.regs[12][10] ),
    .A1(\as1802.regs[13][10] ),
    .A2(\as1802.regs[14][10] ),
    .A3(\as1802.regs[15][10] ),
    .S0(net204),
    .S1(net200),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(_1004_),
    .A1(_1005_),
    .S(net196),
    .X(_1006_));
 sky130_fd_sc_hd__nand2b_1 _4468_ (.A_N(_1006_),
    .B(net194),
    .Y(_1007_));
 sky130_fd_sc_hd__mux4_1 _4469_ (.A0(\as1802.regs[4][10] ),
    .A1(\as1802.regs[5][10] ),
    .A2(\as1802.regs[6][10] ),
    .A3(\as1802.regs[7][10] ),
    .S0(net204),
    .S1(net200),
    .X(_1008_));
 sky130_fd_sc_hd__mux4_1 _4470_ (.A0(\as1802.regs[0][10] ),
    .A1(\as1802.regs[1][10] ),
    .A2(\as1802.regs[2][10] ),
    .A3(\as1802.regs[3][10] ),
    .S0(net205),
    .S1(net201),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(_1009_),
    .A1(_1008_),
    .S(net196),
    .X(_1010_));
 sky130_fd_sc_hd__o21ai_2 _4472_ (.A1(net194),
    .A2(_1010_),
    .B1(_1007_),
    .Y(_1011_));
 sky130_fd_sc_hd__nand2_1 _4473_ (.A(net89),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__or2_1 _4474_ (.A(net89),
    .B(_1011_),
    .X(_1013_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_1012_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a21o_1 _4476_ (.A1(_0829_),
    .A2(_0963_),
    .B1(net89),
    .X(_1015_));
 sky130_fd_sc_hd__or4b_1 _4477_ (.A(_0922_),
    .B(_0964_),
    .C(_0965_),
    .D_N(_0832_),
    .X(_1016_));
 sky130_fd_sc_hd__and2_1 _4478_ (.A(_1015_),
    .B(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__or2_1 _4479_ (.A(_1014_),
    .B(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__a21oi_1 _4480_ (.A1(_1014_),
    .A2(_1017_),
    .B1(_0820_),
    .Y(_1019_));
 sky130_fd_sc_hd__a2bb2o_1 _4481_ (.A1_N(_0462_),
    .A2_N(_0821_),
    .B1(_1018_),
    .B2(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(_1003_),
    .A1(_1020_),
    .S(net81),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_8 _4483_ (.A0(_0983_),
    .A1(_1021_),
    .S(net85),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(net714),
    .A1(_1022_),
    .S(_0705_),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(_0982_),
    .A1(net715),
    .S(_0636_),
    .X(_0030_));
 sky130_fd_sc_hd__or2_1 _4486_ (.A(_0473_),
    .B(_0976_),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _4487_ (.A(_0473_),
    .B(_0976_),
    .Y(_1025_));
 sky130_fd_sc_hd__and2_1 _4488_ (.A(_1024_),
    .B(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__o22a_1 _4489_ (.A1(net130),
    .A2(_0623_),
    .B1(_0979_),
    .B2(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a21o_1 _4490_ (.A1(_0463_),
    .A2(_0473_),
    .B1(_0647_),
    .X(_1028_));
 sky130_fd_sc_hd__o22a_1 _4491_ (.A1(_0624_),
    .A2(_1027_),
    .B1(_1028_),
    .B2(_0474_),
    .X(_1029_));
 sky130_fd_sc_hd__or2_4 _4492_ (.A(net83),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__or3_1 _4493_ (.A(\as1802.regs[2][10] ),
    .B(\as1802.regs[2][11] ),
    .C(_0972_),
    .X(_1031_));
 sky130_fd_sc_hd__o21ai_1 _4494_ (.A1(\as1802.regs[2][10] ),
    .A2(_0972_),
    .B1(net844),
    .Y(_1032_));
 sky130_fd_sc_hd__nand2_1 _4495_ (.A(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__mux4_1 _4496_ (.A0(\as1802.regs[8][11] ),
    .A1(\as1802.regs[9][11] ),
    .A2(\as1802.regs[10][11] ),
    .A3(\as1802.regs[11][11] ),
    .S0(net183),
    .S1(net179),
    .X(_1034_));
 sky130_fd_sc_hd__mux4_1 _4497_ (.A0(\as1802.regs[12][11] ),
    .A1(\as1802.regs[13][11] ),
    .A2(\as1802.regs[14][11] ),
    .A3(\as1802.regs[15][11] ),
    .S0(net183),
    .S1(net179),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(_1034_),
    .A1(_1035_),
    .S(net176),
    .X(_1036_));
 sky130_fd_sc_hd__and2_1 _4499_ (.A(net175),
    .B(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__mux4_1 _4500_ (.A0(\as1802.regs[4][11] ),
    .A1(\as1802.regs[5][11] ),
    .A2(\as1802.regs[6][11] ),
    .A3(\as1802.regs[7][11] ),
    .S0(net183),
    .S1(net179),
    .X(_1038_));
 sky130_fd_sc_hd__mux4_1 _4501_ (.A0(\as1802.regs[0][11] ),
    .A1(\as1802.regs[1][11] ),
    .A2(\as1802.regs[2][11] ),
    .A3(\as1802.regs[3][11] ),
    .S0(net183),
    .S1(net179),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(_1038_),
    .A1(_1039_),
    .S(net113),
    .X(_1040_));
 sky130_fd_sc_hd__a21oi_4 _4503_ (.A1(_3470_),
    .A2(_1040_),
    .B1(_1037_),
    .Y(_1041_));
 sky130_fd_sc_hd__or2_1 _4504_ (.A(_0993_),
    .B(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nor2_1 _4505_ (.A(_0799_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__o21a_1 _4506_ (.A1(_0799_),
    .A2(_0993_),
    .B1(_1041_),
    .X(_1044_));
 sky130_fd_sc_hd__or2_1 _4507_ (.A(_1043_),
    .B(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__nand2_1 _4508_ (.A(_0993_),
    .B(_1041_),
    .Y(_1046_));
 sky130_fd_sc_hd__nand3_1 _4509_ (.A(_0805_),
    .B(_1042_),
    .C(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__o311a_1 _4510_ (.A1(net165),
    .A2(_0573_),
    .A3(_1041_),
    .B1(_1047_),
    .C1(_0675_),
    .X(_1048_));
 sky130_fd_sc_hd__o21a_1 _4511_ (.A1(_0810_),
    .A2(_1045_),
    .B1(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__a211o_1 _4512_ (.A1(net106),
    .A2(_0674_),
    .B1(_1049_),
    .C1(net82),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(_1041_),
    .A1(_1045_),
    .S(net166),
    .X(_1051_));
 sky130_fd_sc_hd__o21ai_1 _4514_ (.A1(_0658_),
    .A2(_1051_),
    .B1(_1050_),
    .Y(_1052_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(net3),
    .A1(_1052_),
    .S(net78),
    .X(_1053_));
 sky130_fd_sc_hd__mux4_1 _4516_ (.A0(\as1802.regs[8][11] ),
    .A1(\as1802.regs[9][11] ),
    .A2(\as1802.regs[10][11] ),
    .A3(\as1802.regs[11][11] ),
    .S0(net204),
    .S1(net200),
    .X(_1054_));
 sky130_fd_sc_hd__mux4_1 _4517_ (.A0(\as1802.regs[12][11] ),
    .A1(\as1802.regs[13][11] ),
    .A2(\as1802.regs[14][11] ),
    .A3(\as1802.regs[15][11] ),
    .S0(net204),
    .S1(net200),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(_1054_),
    .A1(_1055_),
    .S(net196),
    .X(_1056_));
 sky130_fd_sc_hd__mux4_1 _4519_ (.A0(\as1802.regs[4][11] ),
    .A1(\as1802.regs[5][11] ),
    .A2(\as1802.regs[6][11] ),
    .A3(\as1802.regs[7][11] ),
    .S0(net205),
    .S1(net201),
    .X(_1057_));
 sky130_fd_sc_hd__mux4_1 _4520_ (.A0(\as1802.regs[0][11] ),
    .A1(\as1802.regs[1][11] ),
    .A2(\as1802.regs[2][11] ),
    .A3(\as1802.regs[3][11] ),
    .S0(net205),
    .S1(net201),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(_1058_),
    .A1(_1057_),
    .S(net196),
    .X(_1059_));
 sky130_fd_sc_hd__and2b_1 _4522_ (.A_N(net194),
    .B(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__a21oi_2 _4523_ (.A1(net194),
    .A2(_1056_),
    .B1(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__xnor2_1 _4524_ (.A(net90),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_1013_),
    .B(_1018_),
    .Y(_1063_));
 sky130_fd_sc_hd__xnor2_1 _4526_ (.A(_1062_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__mux2_1 _4527_ (.A0(_0473_),
    .A1(_1064_),
    .S(_0821_),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(_1053_),
    .A1(_1065_),
    .S(net81),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_8 _4529_ (.A0(_1033_),
    .A1(_1066_),
    .S(net85),
    .X(_1067_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(net665),
    .A1(_1067_),
    .S(_0705_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(_1030_),
    .A1(net666),
    .S(_0636_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _4532_ (.A(_3608_),
    .B(_1025_),
    .X(_1069_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_3608_),
    .B(_1025_),
    .Y(_1070_));
 sky130_fd_sc_hd__and2_1 _4534_ (.A(_1069_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__o22a_1 _4535_ (.A1(net127),
    .A2(_0623_),
    .B1(_0979_),
    .B2(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__nor2_1 _4536_ (.A(_3608_),
    .B(_0474_),
    .Y(_1073_));
 sky130_fd_sc_hd__o32a_1 _4537_ (.A1(_0475_),
    .A2(_0647_),
    .A3(_1073_),
    .B1(_1072_),
    .B2(_0624_),
    .X(_1074_));
 sky130_fd_sc_hd__or2_4 _4538_ (.A(_0627_),
    .B(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(\as1802.regs[2][12] ),
    .B(_1031_),
    .Y(_1076_));
 sky130_fd_sc_hd__or2_2 _4540_ (.A(\as1802.regs[2][12] ),
    .B(_1031_),
    .X(_1077_));
 sky130_fd_sc_hd__a21oi_1 _4541_ (.A1(_1076_),
    .A2(_1077_),
    .B1(net85),
    .Y(_1078_));
 sky130_fd_sc_hd__mux4_1 _4542_ (.A0(\as1802.regs[8][12] ),
    .A1(\as1802.regs[9][12] ),
    .A2(\as1802.regs[10][12] ),
    .A3(\as1802.regs[11][12] ),
    .S0(net183),
    .S1(net179),
    .X(_1079_));
 sky130_fd_sc_hd__mux4_1 _4543_ (.A0(\as1802.regs[12][12] ),
    .A1(\as1802.regs[13][12] ),
    .A2(\as1802.regs[14][12] ),
    .A3(\as1802.regs[15][12] ),
    .S0(net183),
    .S1(net179),
    .X(_1080_));
 sky130_fd_sc_hd__mux2_1 _4544_ (.A0(_1079_),
    .A1(_1080_),
    .S(net176),
    .X(_1081_));
 sky130_fd_sc_hd__and2_1 _4545_ (.A(net175),
    .B(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__mux4_1 _4546_ (.A0(\as1802.regs[4][12] ),
    .A1(\as1802.regs[5][12] ),
    .A2(\as1802.regs[6][12] ),
    .A3(\as1802.regs[7][12] ),
    .S0(net183),
    .S1(net179),
    .X(_1083_));
 sky130_fd_sc_hd__mux4_1 _4547_ (.A0(\as1802.regs[0][12] ),
    .A1(\as1802.regs[1][12] ),
    .A2(\as1802.regs[2][12] ),
    .A3(\as1802.regs[3][12] ),
    .S0(net183),
    .S1(net179),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _4548_ (.A0(_1083_),
    .A1(_1084_),
    .S(net113),
    .X(_1085_));
 sky130_fd_sc_hd__a21oi_4 _4549_ (.A1(_3470_),
    .A2(_1085_),
    .B1(_1082_),
    .Y(_1086_));
 sky130_fd_sc_hd__inv_2 _4550_ (.A(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__and2b_1 _4551_ (.A_N(_1042_),
    .B(_0809_),
    .X(_1088_));
 sky130_fd_sc_hd__xnor2_1 _4552_ (.A(_1086_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_1043_),
    .B(_1087_),
    .Y(_1090_));
 sky130_fd_sc_hd__xnor2_1 _4554_ (.A(_1043_),
    .B(_1086_),
    .Y(_1091_));
 sky130_fd_sc_hd__mux2_1 _4555_ (.A0(_1091_),
    .A1(_1089_),
    .S(_0810_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _4556_ (.A0(net148),
    .A1(_1092_),
    .S(_0675_),
    .X(_1093_));
 sky130_fd_sc_hd__or2_1 _4557_ (.A(net82),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _4558_ (.A(net165),
    .B(_1086_),
    .Y(_1095_));
 sky130_fd_sc_hd__a211o_1 _4559_ (.A1(net165),
    .A2(_1091_),
    .B1(_1095_),
    .C1(_0658_),
    .X(_1096_));
 sky130_fd_sc_hd__a31o_1 _4560_ (.A1(net4),
    .A2(_0673_),
    .A3(_0675_),
    .B1(net81),
    .X(_1097_));
 sky130_fd_sc_hd__a31o_1 _4561_ (.A1(net78),
    .A2(_1094_),
    .A3(_1096_),
    .B1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__mux4_1 _4562_ (.A0(\as1802.regs[8][12] ),
    .A1(\as1802.regs[9][12] ),
    .A2(\as1802.regs[10][12] ),
    .A3(\as1802.regs[11][12] ),
    .S0(net204),
    .S1(net200),
    .X(_1099_));
 sky130_fd_sc_hd__mux4_1 _4563_ (.A0(\as1802.regs[12][12] ),
    .A1(\as1802.regs[13][12] ),
    .A2(\as1802.regs[14][12] ),
    .A3(\as1802.regs[15][12] ),
    .S0(net204),
    .S1(net200),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _4564_ (.A0(_1099_),
    .A1(_1100_),
    .S(net196),
    .X(_1101_));
 sky130_fd_sc_hd__mux4_1 _4565_ (.A0(\as1802.regs[4][12] ),
    .A1(\as1802.regs[5][12] ),
    .A2(\as1802.regs[6][12] ),
    .A3(\as1802.regs[7][12] ),
    .S0(net205),
    .S1(net201),
    .X(_1102_));
 sky130_fd_sc_hd__mux4_1 _4566_ (.A0(\as1802.regs[0][12] ),
    .A1(\as1802.regs[1][12] ),
    .A2(\as1802.regs[2][12] ),
    .A3(\as1802.regs[3][12] ),
    .S0(net205),
    .S1(net201),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _4567_ (.A0(_1103_),
    .A1(_1102_),
    .S(net196),
    .X(_1104_));
 sky130_fd_sc_hd__and2b_1 _4568_ (.A_N(net194),
    .B(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__a21oi_2 _4569_ (.A1(net194),
    .A2(_1101_),
    .B1(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__and2_1 _4570_ (.A(net90),
    .B(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__nor2_1 _4571_ (.A(net90),
    .B(_1106_),
    .Y(_1108_));
 sky130_fd_sc_hd__nor2_1 _4572_ (.A(_1107_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__inv_2 _4573_ (.A(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__o211a_1 _4574_ (.A1(net90),
    .A2(_1061_),
    .B1(_1015_),
    .C1(_1013_),
    .X(_1111_));
 sky130_fd_sc_hd__o31a_1 _4575_ (.A1(_1014_),
    .A2(_1016_),
    .A3(_1062_),
    .B1(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__and2_1 _4576_ (.A(_1110_),
    .B(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__nor2_1 _4577_ (.A(_1110_),
    .B(_1112_),
    .Y(_1114_));
 sky130_fd_sc_hd__or3_1 _4578_ (.A(_0820_),
    .B(_1113_),
    .C(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__o211ai_1 _4579_ (.A1(_3608_),
    .A2(_0821_),
    .B1(_1115_),
    .C1(net81),
    .Y(_1116_));
 sky130_fd_sc_hd__a31o_4 _4580_ (.A1(net85),
    .A2(_1098_),
    .A3(_1116_),
    .B1(_1078_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(net652),
    .A1(_1117_),
    .S(_0705_),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_1 _4582_ (.A0(_1075_),
    .A1(_1118_),
    .S(_0636_),
    .X(_0032_));
 sky130_fd_sc_hd__nor2_1 _4583_ (.A(_3600_),
    .B(_1069_),
    .Y(_1119_));
 sky130_fd_sc_hd__and2_1 _4584_ (.A(_3600_),
    .B(_1069_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_1 _4585_ (.A(_1119_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__o22a_1 _4586_ (.A1(net125),
    .A2(_0623_),
    .B1(_0979_),
    .B2(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__a21oi_1 _4587_ (.A1(_3608_),
    .A2(_0474_),
    .B1(_3600_),
    .Y(_1123_));
 sky130_fd_sc_hd__o32a_1 _4588_ (.A1(_0476_),
    .A2(_0647_),
    .A3(_1123_),
    .B1(_1122_),
    .B2(_0624_),
    .X(_1124_));
 sky130_fd_sc_hd__or2_4 _4589_ (.A(_0627_),
    .B(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__a21oi_1 _4590_ (.A1(net838),
    .A2(_1077_),
    .B1(net85),
    .Y(_1126_));
 sky130_fd_sc_hd__o21ai_1 _4591_ (.A1(net838),
    .A2(_1077_),
    .B1(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__mux4_1 _4592_ (.A0(\as1802.regs[8][13] ),
    .A1(\as1802.regs[9][13] ),
    .A2(\as1802.regs[10][13] ),
    .A3(\as1802.regs[11][13] ),
    .S0(net183),
    .S1(net179),
    .X(_1128_));
 sky130_fd_sc_hd__mux4_1 _4593_ (.A0(\as1802.regs[12][13] ),
    .A1(\as1802.regs[13][13] ),
    .A2(\as1802.regs[14][13] ),
    .A3(\as1802.regs[15][13] ),
    .S0(net184),
    .S1(net180),
    .X(_1129_));
 sky130_fd_sc_hd__mux2_1 _4594_ (.A0(_1128_),
    .A1(_1129_),
    .S(net176),
    .X(_1130_));
 sky130_fd_sc_hd__and2_1 _4595_ (.A(net175),
    .B(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__mux4_1 _4596_ (.A0(\as1802.regs[4][13] ),
    .A1(\as1802.regs[5][13] ),
    .A2(\as1802.regs[6][13] ),
    .A3(\as1802.regs[7][13] ),
    .S0(net183),
    .S1(net179),
    .X(_1132_));
 sky130_fd_sc_hd__mux4_1 _4597_ (.A0(\as1802.regs[0][13] ),
    .A1(\as1802.regs[1][13] ),
    .A2(\as1802.regs[2][13] ),
    .A3(\as1802.regs[3][13] ),
    .S0(net183),
    .S1(net179),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(_1132_),
    .A1(_1133_),
    .S(net113),
    .X(_1134_));
 sky130_fd_sc_hd__a21oi_4 _4599_ (.A1(_3470_),
    .A2(_1134_),
    .B1(_1131_),
    .Y(_1135_));
 sky130_fd_sc_hd__inv_2 _4600_ (.A(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__or3_2 _4601_ (.A(_1042_),
    .B(_1086_),
    .C(_1135_),
    .X(_1137_));
 sky130_fd_sc_hd__or2_1 _4602_ (.A(_0799_),
    .B(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__a21boi_1 _4603_ (.A1(_1090_),
    .A2(_1135_),
    .B1_N(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__a21oi_1 _4604_ (.A1(_1087_),
    .A2(_1088_),
    .B1(_1136_),
    .Y(_1140_));
 sky130_fd_sc_hd__o21ba_1 _4605_ (.A1(_0806_),
    .A2(_1137_),
    .B1_N(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _4606_ (.A0(_1139_),
    .A1(_1141_),
    .S(_0810_),
    .X(_1142_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(_3476_),
    .B(_0674_),
    .Y(_1143_));
 sky130_fd_sc_hd__o211a_1 _4608_ (.A1(_0674_),
    .A2(_1142_),
    .B1(_1143_),
    .C1(_0658_),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _4609_ (.A0(_1136_),
    .A1(_1139_),
    .S(net165),
    .X(_1145_));
 sky130_fd_sc_hd__a21o_1 _4610_ (.A1(net82),
    .A2(_1145_),
    .B1(_0653_),
    .X(_1146_));
 sky130_fd_sc_hd__o22a_1 _4611_ (.A1(_0654_),
    .A2(_1139_),
    .B1(_1144_),
    .B2(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__or2_1 _4612_ (.A(net5),
    .B(_0677_),
    .X(_1148_));
 sky130_fd_sc_hd__o211a_1 _4613_ (.A1(_0676_),
    .A2(_1147_),
    .B1(_1148_),
    .C1(net80),
    .X(_1149_));
 sky130_fd_sc_hd__mux4_1 _4614_ (.A0(\as1802.regs[8][13] ),
    .A1(\as1802.regs[9][13] ),
    .A2(\as1802.regs[10][13] ),
    .A3(\as1802.regs[11][13] ),
    .S0(net204),
    .S1(net200),
    .X(_1150_));
 sky130_fd_sc_hd__mux4_1 _4615_ (.A0(\as1802.regs[12][13] ),
    .A1(\as1802.regs[13][13] ),
    .A2(\as1802.regs[14][13] ),
    .A3(\as1802.regs[15][13] ),
    .S0(net205),
    .S1(net201),
    .X(_1151_));
 sky130_fd_sc_hd__mux2_1 _4616_ (.A0(_1150_),
    .A1(_1151_),
    .S(net196),
    .X(_1152_));
 sky130_fd_sc_hd__mux4_1 _4617_ (.A0(\as1802.regs[4][13] ),
    .A1(\as1802.regs[5][13] ),
    .A2(\as1802.regs[6][13] ),
    .A3(\as1802.regs[7][13] ),
    .S0(net205),
    .S1(net201),
    .X(_1153_));
 sky130_fd_sc_hd__mux4_1 _4618_ (.A0(\as1802.regs[0][13] ),
    .A1(\as1802.regs[1][13] ),
    .A2(\as1802.regs[2][13] ),
    .A3(\as1802.regs[3][13] ),
    .S0(net205),
    .S1(net201),
    .X(_1154_));
 sky130_fd_sc_hd__mux2_1 _4619_ (.A0(_1154_),
    .A1(_1153_),
    .S(net196),
    .X(_1155_));
 sky130_fd_sc_hd__and2b_1 _4620_ (.A_N(net194),
    .B(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a21oi_2 _4621_ (.A1(net194),
    .A2(_1152_),
    .B1(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__and2_1 _4622_ (.A(net90),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__nor2_1 _4623_ (.A(net90),
    .B(_1157_),
    .Y(_1159_));
 sky130_fd_sc_hd__nor2_1 _4624_ (.A(_1158_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__or3_1 _4625_ (.A(_1108_),
    .B(_1114_),
    .C(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__o21ai_1 _4626_ (.A1(_1108_),
    .A2(_1114_),
    .B1(_1160_),
    .Y(_1162_));
 sky130_fd_sc_hd__a21oi_1 _4627_ (.A1(_1161_),
    .A2(_1162_),
    .B1(_0820_),
    .Y(_1163_));
 sky130_fd_sc_hd__a211oi_1 _4628_ (.A1(_3600_),
    .A2(_0820_),
    .B1(_1163_),
    .C1(_0685_),
    .Y(_1164_));
 sky130_fd_sc_hd__o31a_4 _4629_ (.A1(_0687_),
    .A2(_1149_),
    .A3(_1164_),
    .B1(_1127_),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(net650),
    .A1(_1165_),
    .S(_0705_),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(_1125_),
    .A1(net651),
    .S(_0636_),
    .X(_0033_));
 sky130_fd_sc_hd__or3_1 _4632_ (.A(_3592_),
    .B(_3600_),
    .C(_1069_),
    .X(_1167_));
 sky130_fd_sc_hd__xnor2_1 _4633_ (.A(_3592_),
    .B(_1119_),
    .Y(_1168_));
 sky130_fd_sc_hd__o22a_1 _4634_ (.A1(net122),
    .A2(_0623_),
    .B1(_0979_),
    .B2(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__o21a_1 _4635_ (.A1(_3592_),
    .A2(_0476_),
    .B1(_0648_),
    .X(_1170_));
 sky130_fd_sc_hd__o2bb2a_1 _4636_ (.A1_N(_0477_),
    .A2_N(_1170_),
    .B1(_1169_),
    .B2(_0624_),
    .X(_1171_));
 sky130_fd_sc_hd__or2_4 _4637_ (.A(_0627_),
    .B(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__or3_1 _4638_ (.A(\as1802.regs[2][13] ),
    .B(\as1802.regs[2][14] ),
    .C(_1077_),
    .X(_1173_));
 sky130_fd_sc_hd__o21ai_1 _4639_ (.A1(net886),
    .A2(_1077_),
    .B1(\as1802.regs[2][14] ),
    .Y(_1174_));
 sky130_fd_sc_hd__a21oi_1 _4640_ (.A1(_1173_),
    .A2(_1174_),
    .B1(net85),
    .Y(_1175_));
 sky130_fd_sc_hd__mux4_1 _4641_ (.A0(\as1802.regs[8][14] ),
    .A1(\as1802.regs[9][14] ),
    .A2(\as1802.regs[10][14] ),
    .A3(\as1802.regs[11][14] ),
    .S0(net183),
    .S1(net179),
    .X(_1176_));
 sky130_fd_sc_hd__mux4_1 _4642_ (.A0(\as1802.regs[12][14] ),
    .A1(\as1802.regs[13][14] ),
    .A2(\as1802.regs[14][14] ),
    .A3(\as1802.regs[15][14] ),
    .S0(net184),
    .S1(net180),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_1 _4643_ (.A0(_1176_),
    .A1(_1177_),
    .S(net176),
    .X(_1178_));
 sky130_fd_sc_hd__and2_1 _4644_ (.A(net175),
    .B(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__mux4_1 _4645_ (.A0(\as1802.regs[4][14] ),
    .A1(\as1802.regs[5][14] ),
    .A2(\as1802.regs[6][14] ),
    .A3(\as1802.regs[7][14] ),
    .S0(net183),
    .S1(net179),
    .X(_1180_));
 sky130_fd_sc_hd__mux4_1 _4646_ (.A0(\as1802.regs[0][14] ),
    .A1(\as1802.regs[1][14] ),
    .A2(\as1802.regs[2][14] ),
    .A3(\as1802.regs[3][14] ),
    .S0(net183),
    .S1(net179),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_1 _4647_ (.A0(_1180_),
    .A1(_1181_),
    .S(net113),
    .X(_1182_));
 sky130_fd_sc_hd__a21oi_4 _4648_ (.A1(_3470_),
    .A2(_1182_),
    .B1(_1179_),
    .Y(_1183_));
 sky130_fd_sc_hd__inv_2 _4649_ (.A(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__or2_1 _4650_ (.A(_1137_),
    .B(_1183_),
    .X(_1185_));
 sky130_fd_sc_hd__nor2_1 _4651_ (.A(_0799_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a21oi_1 _4652_ (.A1(_1138_),
    .A2(_1183_),
    .B1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__or2_1 _4653_ (.A(net165),
    .B(_1183_),
    .X(_1188_));
 sky130_fd_sc_hd__inv_2 _4654_ (.A(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4655_ (.A(_1137_),
    .B(_1183_),
    .Y(_1190_));
 sky130_fd_sc_hd__a32o_1 _4656_ (.A1(_0805_),
    .A2(_1185_),
    .A3(_1190_),
    .B1(_1189_),
    .B2(_0572_),
    .X(_1191_));
 sky130_fd_sc_hd__a21oi_1 _4657_ (.A1(_0807_),
    .A2(_1187_),
    .B1(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__nor2_1 _4658_ (.A(_0674_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__a211o_1 _4659_ (.A1(net142),
    .A2(_0674_),
    .B1(_1193_),
    .C1(_0657_),
    .X(_1194_));
 sky130_fd_sc_hd__a211o_1 _4660_ (.A1(net165),
    .A2(_1187_),
    .B1(_1189_),
    .C1(_0658_),
    .X(_1195_));
 sky130_fd_sc_hd__a21o_1 _4661_ (.A1(_1194_),
    .A2(_1195_),
    .B1(_0653_),
    .X(_1196_));
 sky130_fd_sc_hd__o21a_1 _4662_ (.A1(_0654_),
    .A2(_1187_),
    .B1(net78),
    .X(_1197_));
 sky130_fd_sc_hd__a221o_1 _4663_ (.A1(net6),
    .A2(_0676_),
    .B1(_1196_),
    .B2(_1197_),
    .C1(net81),
    .X(_1198_));
 sky130_fd_sc_hd__mux4_1 _4664_ (.A0(\as1802.regs[8][14] ),
    .A1(\as1802.regs[9][14] ),
    .A2(\as1802.regs[10][14] ),
    .A3(\as1802.regs[11][14] ),
    .S0(net204),
    .S1(net200),
    .X(_1199_));
 sky130_fd_sc_hd__mux4_1 _4665_ (.A0(\as1802.regs[12][14] ),
    .A1(\as1802.regs[13][14] ),
    .A2(\as1802.regs[14][14] ),
    .A3(\as1802.regs[15][14] ),
    .S0(_0004_),
    .S1(_0005_),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _4666_ (.A0(_1199_),
    .A1(_1200_),
    .S(net196),
    .X(_1201_));
 sky130_fd_sc_hd__nand2b_1 _4667_ (.A_N(_1201_),
    .B(net194),
    .Y(_1202_));
 sky130_fd_sc_hd__mux4_1 _4668_ (.A0(\as1802.regs[4][14] ),
    .A1(\as1802.regs[5][14] ),
    .A2(\as1802.regs[6][14] ),
    .A3(\as1802.regs[7][14] ),
    .S0(net205),
    .S1(net201),
    .X(_1203_));
 sky130_fd_sc_hd__mux4_1 _4669_ (.A0(\as1802.regs[0][14] ),
    .A1(\as1802.regs[1][14] ),
    .A2(\as1802.regs[2][14] ),
    .A3(\as1802.regs[3][14] ),
    .S0(net205),
    .S1(net201),
    .X(_1204_));
 sky130_fd_sc_hd__mux2_1 _4670_ (.A0(_1204_),
    .A1(_1203_),
    .S(net196),
    .X(_1205_));
 sky130_fd_sc_hd__o21ai_2 _4671_ (.A1(net194),
    .A2(_1205_),
    .B1(_1202_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2b_1 _4672_ (.A_N(_1206_),
    .B(net90),
    .Y(_1207_));
 sky130_fd_sc_hd__nand2b_1 _4673_ (.A_N(net90),
    .B(_1206_),
    .Y(_1208_));
 sky130_fd_sc_hd__and2_1 _4674_ (.A(_1207_),
    .B(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__a211o_1 _4675_ (.A1(_1114_),
    .A2(_1160_),
    .B1(_1159_),
    .C1(_1108_),
    .X(_1210_));
 sky130_fd_sc_hd__xnor2_1 _4676_ (.A(_1209_),
    .B(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__nor2_1 _4677_ (.A(_3592_),
    .B(_0821_),
    .Y(_1212_));
 sky130_fd_sc_hd__a211o_1 _4678_ (.A1(_0821_),
    .A2(_1211_),
    .B1(_1212_),
    .C1(_0685_),
    .X(_1213_));
 sky130_fd_sc_hd__a31o_4 _4679_ (.A1(net85),
    .A2(_1198_),
    .A3(_1213_),
    .B1(_1175_),
    .X(_1214_));
 sky130_fd_sc_hd__mux2_1 _4680_ (.A0(net689),
    .A1(_1214_),
    .S(_0705_),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _4681_ (.A0(_1172_),
    .A1(_1215_),
    .S(_0636_),
    .X(_0034_));
 sky130_fd_sc_hd__xor2_1 _4682_ (.A(_0485_),
    .B(_1167_),
    .X(_1216_));
 sky130_fd_sc_hd__o22a_1 _4683_ (.A1(net120),
    .A2(_0623_),
    .B1(_0979_),
    .B2(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__o2bb2a_1 _4684_ (.A1_N(_0486_),
    .A2_N(_0648_),
    .B1(_1217_),
    .B2(_0624_),
    .X(_1218_));
 sky130_fd_sc_hd__or2_4 _4685_ (.A(_0627_),
    .B(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__mux4_1 _4686_ (.A0(\as1802.regs[8][15] ),
    .A1(\as1802.regs[9][15] ),
    .A2(\as1802.regs[10][15] ),
    .A3(\as1802.regs[11][15] ),
    .S0(net184),
    .S1(net180),
    .X(_1220_));
 sky130_fd_sc_hd__mux4_1 _4687_ (.A0(\as1802.regs[12][15] ),
    .A1(\as1802.regs[13][15] ),
    .A2(\as1802.regs[14][15] ),
    .A3(\as1802.regs[15][15] ),
    .S0(_0008_),
    .S1(_0009_),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _4688_ (.A0(_1220_),
    .A1(_1221_),
    .S(net176),
    .X(_1222_));
 sky130_fd_sc_hd__and2_1 _4689_ (.A(net175),
    .B(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__mux4_1 _4690_ (.A0(\as1802.regs[4][15] ),
    .A1(\as1802.regs[5][15] ),
    .A2(\as1802.regs[6][15] ),
    .A3(\as1802.regs[7][15] ),
    .S0(net183),
    .S1(net179),
    .X(_1224_));
 sky130_fd_sc_hd__mux4_1 _4691_ (.A0(\as1802.regs[0][15] ),
    .A1(\as1802.regs[1][15] ),
    .A2(\as1802.regs[2][15] ),
    .A3(\as1802.regs[3][15] ),
    .S0(net183),
    .S1(net179),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _4692_ (.A0(_1224_),
    .A1(_1225_),
    .S(net113),
    .X(_1226_));
 sky130_fd_sc_hd__a21oi_2 _4693_ (.A1(_3470_),
    .A2(_1226_),
    .B1(_1223_),
    .Y(_1227_));
 sky130_fd_sc_hd__inv_2 _4694_ (.A(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__xnor2_1 _4695_ (.A(_1186_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__a21o_1 _4696_ (.A1(net118),
    .A2(_1227_),
    .B1(_0658_),
    .X(_1230_));
 sky130_fd_sc_hd__a21o_1 _4697_ (.A1(net166),
    .A2(_1229_),
    .B1(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__or3_1 _4698_ (.A(_0806_),
    .B(_1137_),
    .C(_1183_),
    .X(_1232_));
 sky130_fd_sc_hd__xnor2_1 _4699_ (.A(_1228_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__nor2_1 _4700_ (.A(net139),
    .B(_0675_),
    .Y(_1234_));
 sky130_fd_sc_hd__or4_1 _4701_ (.A(net82),
    .B(_0810_),
    .C(_1229_),
    .D(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a21oi_1 _4702_ (.A1(_0810_),
    .A2(_1233_),
    .B1(_0674_),
    .Y(_1236_));
 sky130_fd_sc_hd__o211a_1 _4703_ (.A1(_1234_),
    .A2(_1236_),
    .B1(net78),
    .C1(_1231_),
    .X(_1237_));
 sky130_fd_sc_hd__a221o_1 _4704_ (.A1(_3479_),
    .A2(_0676_),
    .B1(_1235_),
    .B2(_1237_),
    .C1(net81),
    .X(_1238_));
 sky130_fd_sc_hd__mux4_1 _4705_ (.A0(\as1802.regs[8][15] ),
    .A1(\as1802.regs[9][15] ),
    .A2(\as1802.regs[10][15] ),
    .A3(\as1802.regs[11][15] ),
    .S0(_0004_),
    .S1(_0005_),
    .X(_1239_));
 sky130_fd_sc_hd__mux4_1 _4706_ (.A0(\as1802.regs[12][15] ),
    .A1(\as1802.regs[13][15] ),
    .A2(\as1802.regs[14][15] ),
    .A3(\as1802.regs[15][15] ),
    .S0(net204),
    .S1(net200),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(_1239_),
    .A1(_1240_),
    .S(net196),
    .X(_1241_));
 sky130_fd_sc_hd__mux4_1 _4708_ (.A0(\as1802.regs[4][15] ),
    .A1(\as1802.regs[5][15] ),
    .A2(\as1802.regs[6][15] ),
    .A3(\as1802.regs[7][15] ),
    .S0(net205),
    .S1(net201),
    .X(_1242_));
 sky130_fd_sc_hd__mux4_1 _4709_ (.A0(\as1802.regs[0][15] ),
    .A1(\as1802.regs[1][15] ),
    .A2(\as1802.regs[2][15] ),
    .A3(\as1802.regs[3][15] ),
    .S0(net205),
    .S1(net201),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _4710_ (.A0(_1243_),
    .A1(_1242_),
    .S(net196),
    .X(_1244_));
 sky130_fd_sc_hd__and2b_1 _4711_ (.A_N(net195),
    .B(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__a21oi_2 _4712_ (.A1(_0007_),
    .A2(_1241_),
    .B1(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__mux2_1 _4713_ (.A0(_1208_),
    .A1(_1207_),
    .S(_1210_),
    .X(_1247_));
 sky130_fd_sc_hd__xnor2_1 _4714_ (.A(_1246_),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__mux2_1 _4715_ (.A0(_0485_),
    .A1(_1248_),
    .S(_0821_),
    .X(_1249_));
 sky130_fd_sc_hd__a21oi_1 _4716_ (.A1(\as1802.regs[2][15] ),
    .A2(_1173_),
    .B1(net85),
    .Y(_1250_));
 sky130_fd_sc_hd__o21a_1 _4717_ (.A1(\as1802.regs[2][15] ),
    .A2(_1173_),
    .B1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__o211a_2 _4718_ (.A1(_0685_),
    .A2(_1249_),
    .B1(_1238_),
    .C1(net85),
    .X(_1252_));
 sky130_fd_sc_hd__nor2_8 _4719_ (.A(_1251_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__mux2_1 _4720_ (.A0(net800),
    .A1(_1253_),
    .S(_0705_),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(_1219_),
    .A1(_1254_),
    .S(_0636_),
    .X(_0035_));
 sky130_fd_sc_hd__a21boi_1 _4722_ (.A1(_3480_),
    .A2(_3559_),
    .B1_N(_3560_),
    .Y(_0036_));
 sky130_fd_sc_hd__nor2_1 _4723_ (.A(net103),
    .B(_3540_),
    .Y(_1255_));
 sky130_fd_sc_hd__mux2_1 _4724_ (.A0(_1255_),
    .A1(net817),
    .S(_3559_),
    .X(_0037_));
 sky130_fd_sc_hd__and2b_2 _4725_ (.A_N(_0629_),
    .B(_0628_),
    .X(_1256_));
 sky130_fd_sc_hd__and2b_2 _4726_ (.A_N(_0632_),
    .B(_0631_),
    .X(_1257_));
 sky130_fd_sc_hd__and3_4 _4727_ (.A(_0635_),
    .B(_1256_),
    .C(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__and3_2 _4728_ (.A(net84),
    .B(_0689_),
    .C(_0693_),
    .X(_1259_));
 sky130_fd_sc_hd__nor2_4 _4729_ (.A(_0698_),
    .B(_0701_),
    .Y(_1260_));
 sky130_fd_sc_hd__and3_4 _4730_ (.A(_0704_),
    .B(_1259_),
    .C(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__mux2_1 _4731_ (.A0(net482),
    .A1(_0926_),
    .S(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__mux2_1 _4732_ (.A0(net483),
    .A1(_0652_),
    .S(_1258_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4733_ (.A0(net675),
    .A1(_0974_),
    .S(_1261_),
    .X(_1263_));
 sky130_fd_sc_hd__mux2_1 _4734_ (.A0(_1263_),
    .A1(_0934_),
    .S(_1258_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4735_ (.A0(net589),
    .A1(_1022_),
    .S(_1261_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_1 _4736_ (.A0(net590),
    .A1(_0982_),
    .S(_1258_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4737_ (.A0(net562),
    .A1(_1067_),
    .S(_1261_),
    .X(_1265_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(net563),
    .A1(_1030_),
    .S(_1258_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(net436),
    .A1(_1117_),
    .S(_1261_),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _4740_ (.A0(_1266_),
    .A1(_1075_),
    .S(_1258_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(net736),
    .A1(_1165_),
    .S(_1261_),
    .X(_1267_));
 sky130_fd_sc_hd__mux2_1 _4742_ (.A0(net737),
    .A1(_1125_),
    .S(_1258_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4743_ (.A0(net421),
    .A1(_1214_),
    .S(_1261_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(_1268_),
    .A1(_1172_),
    .S(_1258_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4745_ (.A0(net433),
    .A1(_1253_),
    .S(_1261_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _4746_ (.A0(_1269_),
    .A1(_1219_),
    .S(_1258_),
    .X(_0045_));
 sky130_fd_sc_hd__nor2_2 _4747_ (.A(_0628_),
    .B(_0629_),
    .Y(_1270_));
 sky130_fd_sc_hd__nor2_4 _4748_ (.A(_0631_),
    .B(_0632_),
    .Y(_1271_));
 sky130_fd_sc_hd__and3_4 _4749_ (.A(_0635_),
    .B(_1270_),
    .C(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__and2_2 _4750_ (.A(_0690_),
    .B(_0693_),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_4 _4751_ (.A(_0697_),
    .B(_0701_),
    .Y(_1274_));
 sky130_fd_sc_hd__and3_4 _4752_ (.A(_0704_),
    .B(_1273_),
    .C(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _4753_ (.A0(net570),
    .A1(_0926_),
    .S(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _4754_ (.A0(net571),
    .A1(_0652_),
    .S(_1272_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4755_ (.A0(net446),
    .A1(_0974_),
    .S(_1275_),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_1 _4756_ (.A0(_1277_),
    .A1(_0934_),
    .S(_1272_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4757_ (.A0(net525),
    .A1(_1022_),
    .S(_1275_),
    .X(_1278_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(net526),
    .A1(_0982_),
    .S(_1272_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4759_ (.A0(net687),
    .A1(_1067_),
    .S(_1275_),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _4760_ (.A0(net688),
    .A1(_1030_),
    .S(_1272_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4761_ (.A0(net663),
    .A1(_1117_),
    .S(_1275_),
    .X(_1280_));
 sky130_fd_sc_hd__mux2_1 _4762_ (.A0(_1280_),
    .A1(_1075_),
    .S(_1272_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4763_ (.A0(net566),
    .A1(_1165_),
    .S(_1275_),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _4764_ (.A0(net567),
    .A1(_1125_),
    .S(_1272_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(net581),
    .A1(_1214_),
    .S(_1275_),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(_1282_),
    .A1(_1172_),
    .S(_1272_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4767_ (.A0(net713),
    .A1(_1253_),
    .S(_1275_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _4768_ (.A0(_1283_),
    .A1(_1219_),
    .S(_1272_),
    .X(_0053_));
 sky130_fd_sc_hd__and3_4 _4769_ (.A(_0635_),
    .B(_1256_),
    .C(_1271_),
    .X(_1284_));
 sky130_fd_sc_hd__and3_4 _4770_ (.A(_0704_),
    .B(_1259_),
    .C(_1274_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _4771_ (.A0(net604),
    .A1(_0926_),
    .S(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _4772_ (.A0(net605),
    .A1(_0652_),
    .S(_1284_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _4773_ (.A0(net603),
    .A1(_0974_),
    .S(_1285_),
    .X(_1287_));
 sky130_fd_sc_hd__mux2_1 _4774_ (.A0(_1287_),
    .A1(_0934_),
    .S(_1284_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _4775_ (.A0(net443),
    .A1(_1022_),
    .S(_1285_),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_1 _4776_ (.A0(net444),
    .A1(_0982_),
    .S(_1284_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4777_ (.A0(net480),
    .A1(_1067_),
    .S(_1285_),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(net481),
    .A1(_1030_),
    .S(_1284_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _4779_ (.A0(net767),
    .A1(_1117_),
    .S(_1285_),
    .X(_1290_));
 sky130_fd_sc_hd__mux2_1 _4780_ (.A0(_1290_),
    .A1(_1075_),
    .S(_1284_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _4781_ (.A0(net531),
    .A1(_1165_),
    .S(_1285_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _4782_ (.A0(net532),
    .A1(_1125_),
    .S(_1284_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4783_ (.A0(net693),
    .A1(_1214_),
    .S(_1285_),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _4784_ (.A0(_1292_),
    .A1(_1172_),
    .S(_1284_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4785_ (.A0(net597),
    .A1(_1253_),
    .S(_1285_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _4786_ (.A0(_1293_),
    .A1(_1219_),
    .S(_1284_),
    .X(_0061_));
 sky130_fd_sc_hd__and2b_2 _4787_ (.A_N(_0628_),
    .B(_0629_),
    .X(_1294_));
 sky130_fd_sc_hd__or3b_4 _4788_ (.A(_0633_),
    .B(_0634_),
    .C_N(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__and3_2 _4789_ (.A(net84),
    .B(_0690_),
    .C(_0692_),
    .X(_1296_));
 sky130_fd_sc_hd__and3_4 _4790_ (.A(_0702_),
    .B(_0704_),
    .C(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_1 _4791_ (.A0(net643),
    .A1(_0926_),
    .S(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__mux2_1 _4792_ (.A0(_0652_),
    .A1(net644),
    .S(_1295_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _4793_ (.A0(net546),
    .A1(_0974_),
    .S(_1297_),
    .X(_1299_));
 sky130_fd_sc_hd__mux2_1 _4794_ (.A0(_0934_),
    .A1(_1299_),
    .S(_1295_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4795_ (.A0(net690),
    .A1(_1022_),
    .S(_1297_),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _4796_ (.A0(_0982_),
    .A1(net691),
    .S(_1295_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _4797_ (.A0(net560),
    .A1(_1067_),
    .S(_1297_),
    .X(_1301_));
 sky130_fd_sc_hd__mux2_1 _4798_ (.A0(_1030_),
    .A1(net561),
    .S(_1295_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4799_ (.A0(net632),
    .A1(_1117_),
    .S(_1297_),
    .X(_1302_));
 sky130_fd_sc_hd__mux2_1 _4800_ (.A0(_1075_),
    .A1(_1302_),
    .S(_1295_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _4801_ (.A0(net610),
    .A1(_1165_),
    .S(_1297_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(_1125_),
    .A1(net611),
    .S(_1295_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(net624),
    .A1(_1214_),
    .S(_1297_),
    .X(_1304_));
 sky130_fd_sc_hd__mux2_1 _4804_ (.A0(_1172_),
    .A1(_1304_),
    .S(_1295_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4805_ (.A0(net674),
    .A1(_1253_),
    .S(_1297_),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(_1219_),
    .A1(_1305_),
    .S(_1295_),
    .X(_0069_));
 sky130_fd_sc_hd__and3_4 _4807_ (.A(_0635_),
    .B(_1257_),
    .C(_1294_),
    .X(_1306_));
 sky130_fd_sc_hd__and3_4 _4808_ (.A(_0704_),
    .B(_1260_),
    .C(_1296_),
    .X(_1307_));
 sky130_fd_sc_hd__mux2_1 _4809_ (.A0(net434),
    .A1(_0926_),
    .S(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(net435),
    .A1(_0652_),
    .S(_1306_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4811_ (.A0(net442),
    .A1(_0974_),
    .S(_1307_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(_1309_),
    .A1(_0934_),
    .S(_1306_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4813_ (.A0(net498),
    .A1(_1022_),
    .S(_1307_),
    .X(_1310_));
 sky130_fd_sc_hd__mux2_1 _4814_ (.A0(net499),
    .A1(_0982_),
    .S(_1306_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4815_ (.A0(net400),
    .A1(_1067_),
    .S(_1307_),
    .X(_1311_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(net401),
    .A1(_1030_),
    .S(_1306_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(net429),
    .A1(_1117_),
    .S(_1307_),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_1 _4818_ (.A0(_1312_),
    .A1(_1075_),
    .S(_1306_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4819_ (.A0(net464),
    .A1(_1165_),
    .S(_1307_),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(net465),
    .A1(_1125_),
    .S(_1306_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _4821_ (.A0(net459),
    .A1(_1214_),
    .S(_1307_),
    .X(_1314_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_1314_),
    .A1(_1172_),
    .S(_1306_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(net704),
    .A1(_1253_),
    .S(_1307_),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _4824_ (.A0(_1315_),
    .A1(_1219_),
    .S(_1306_),
    .X(_0077_));
 sky130_fd_sc_hd__and2b_2 _4825_ (.A_N(_0631_),
    .B(_0632_),
    .X(_1316_));
 sky130_fd_sc_hd__and3_4 _4826_ (.A(_0635_),
    .B(_1294_),
    .C(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__and2_2 _4827_ (.A(_0698_),
    .B(_0701_),
    .X(_1318_));
 sky130_fd_sc_hd__and3_4 _4828_ (.A(_0704_),
    .B(_1296_),
    .C(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _4829_ (.A0(net796),
    .A1(_0926_),
    .S(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__mux2_1 _4830_ (.A0(net797),
    .A1(_0652_),
    .S(_1317_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4831_ (.A0(net439),
    .A1(_0974_),
    .S(_1319_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _4832_ (.A0(_1321_),
    .A1(_0934_),
    .S(_1317_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4833_ (.A0(net490),
    .A1(_1022_),
    .S(_1319_),
    .X(_1322_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(net491),
    .A1(_0982_),
    .S(_1317_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(net412),
    .A1(_1067_),
    .S(_1319_),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_1 _4836_ (.A0(net413),
    .A1(_1030_),
    .S(_1317_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _4837_ (.A0(net411),
    .A1(_1117_),
    .S(_1319_),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(_1324_),
    .A1(_1075_),
    .S(_1317_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4839_ (.A0(net711),
    .A1(_1165_),
    .S(_1319_),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _4840_ (.A0(net712),
    .A1(_1125_),
    .S(_1317_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(net430),
    .A1(_1214_),
    .S(_1319_),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_1 _4842_ (.A0(_1326_),
    .A1(_1172_),
    .S(_1317_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4843_ (.A0(net788),
    .A1(_1253_),
    .S(_1319_),
    .X(_1327_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(_1327_),
    .A1(_1219_),
    .S(_1317_),
    .X(_0085_));
 sky130_fd_sc_hd__and3_2 _4845_ (.A(net211),
    .B(_0622_),
    .C(_0626_),
    .X(_1328_));
 sky130_fd_sc_hd__nand3_4 _4846_ (.A(net211),
    .B(_0622_),
    .C(_0626_),
    .Y(_1329_));
 sky130_fd_sc_hd__and3_4 _4847_ (.A(_1257_),
    .B(_1294_),
    .C(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(net135),
    .A1(_0420_),
    .S(_0622_),
    .X(_1331_));
 sky130_fd_sc_hd__or2_4 _4849_ (.A(net83),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__nand2_8 _4850_ (.A(_0673_),
    .B(_0703_),
    .Y(_1333_));
 sky130_fd_sc_hd__and3_4 _4851_ (.A(_1260_),
    .B(_1296_),
    .C(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__or2_2 _4852_ (.A(net118),
    .B(_0799_),
    .X(_1335_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(net118),
    .B(_0799_),
    .Y(_1336_));
 sky130_fd_sc_hd__a21o_1 _4854_ (.A1(_1335_),
    .A2(_1336_),
    .B1(_0658_),
    .X(_1337_));
 sky130_fd_sc_hd__o21ai_1 _4855_ (.A1(_0799_),
    .A2(_0804_),
    .B1(_0663_),
    .Y(_1338_));
 sky130_fd_sc_hd__o211ai_1 _4856_ (.A1(net111),
    .A2(_0663_),
    .B1(_0806_),
    .C1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__o211a_1 _4857_ (.A1(_0800_),
    .A2(_0807_),
    .B1(_1339_),
    .C1(_0662_),
    .X(_1340_));
 sky130_fd_sc_hd__a211o_1 _4858_ (.A1(net160),
    .A2(_0661_),
    .B1(_1340_),
    .C1(net82),
    .X(_1341_));
 sky130_fd_sc_hd__a21o_1 _4859_ (.A1(_1337_),
    .A2(_1341_),
    .B1(_0676_),
    .X(_1342_));
 sky130_fd_sc_hd__o211a_1 _4860_ (.A1(net1),
    .A2(net78),
    .B1(net80),
    .C1(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__or2_1 _4861_ (.A(_0820_),
    .B(_0889_),
    .X(_1344_));
 sky130_fd_sc_hd__nand2_1 _4862_ (.A(_0420_),
    .B(_0820_),
    .Y(_1345_));
 sky130_fd_sc_hd__a31o_1 _4863_ (.A1(net81),
    .A2(_1344_),
    .A3(_1345_),
    .B1(_0687_),
    .X(_1346_));
 sky130_fd_sc_hd__o22a_4 _4864_ (.A1(_3465_),
    .A2(net84),
    .B1(_1343_),
    .B2(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__mux2_1 _4865_ (.A0(net389),
    .A1(_1347_),
    .S(_1334_),
    .X(_1348_));
 sky130_fd_sc_hd__mux2_1 _4866_ (.A0(net390),
    .A1(_1332_),
    .S(_1330_),
    .X(_0086_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_0429_),
    .B(_0637_),
    .Y(_1349_));
 sky130_fd_sc_hd__xnor2_1 _4868_ (.A(_0646_),
    .B(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(_3437_),
    .A1(_1350_),
    .S(_0622_),
    .X(_1351_));
 sky130_fd_sc_hd__a21oi_1 _4870_ (.A1(_0624_),
    .A2(_1351_),
    .B1(net83),
    .Y(_1352_));
 sky130_fd_sc_hd__o21ai_4 _4871_ (.A1(_0624_),
    .A2(_1351_),
    .B1(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__xnor2_1 _4872_ (.A(\as1802.regs[2][0] ),
    .B(net836),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2_1 _4873_ (.A(_0729_),
    .B(_0799_),
    .Y(_1355_));
 sky130_fd_sc_hd__nor2_1 _4874_ (.A(_0730_),
    .B(_0800_),
    .Y(_1356_));
 sky130_fd_sc_hd__nor2_1 _4875_ (.A(_1355_),
    .B(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__or3b_4 _4876_ (.A(_0572_),
    .B(_0805_),
    .C_N(_0663_),
    .X(_1358_));
 sky130_fd_sc_hd__a22oi_2 _4877_ (.A1(_0729_),
    .A2(_1335_),
    .B1(_1355_),
    .B2(net166),
    .Y(_1359_));
 sky130_fd_sc_hd__o22a_1 _4878_ (.A1(net157),
    .A2(_0663_),
    .B1(_1359_),
    .B2(_0573_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _4879_ (.A0(_1360_),
    .A1(_0729_),
    .S(_0809_),
    .X(_1361_));
 sky130_fd_sc_hd__o211a_1 _4880_ (.A1(_1357_),
    .A2(_1358_),
    .B1(_1361_),
    .C1(_0662_),
    .X(_1362_));
 sky130_fd_sc_hd__a21o_1 _4881_ (.A1(net157),
    .A2(_0661_),
    .B1(net82),
    .X(_1363_));
 sky130_fd_sc_hd__o22a_1 _4882_ (.A1(_0658_),
    .A2(_1359_),
    .B1(_1362_),
    .B2(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(net12),
    .A1(_1364_),
    .S(net78),
    .X(_1365_));
 sky130_fd_sc_hd__a21o_1 _4884_ (.A1(_0881_),
    .A2(_0889_),
    .B1(_0820_),
    .X(_1366_));
 sky130_fd_sc_hd__o221a_1 _4885_ (.A1(_0428_),
    .A2(_0821_),
    .B1(_0890_),
    .B2(_1366_),
    .C1(net81),
    .X(_1367_));
 sky130_fd_sc_hd__o21ba_1 _4886_ (.A1(net81),
    .A2(_1365_),
    .B1_N(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_8 _4887_ (.A0(_1354_),
    .A1(_1368_),
    .S(net84),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_1 _4888_ (.A0(net547),
    .A1(_1369_),
    .S(_1334_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _4889_ (.A0(net548),
    .A1(_1353_),
    .S(_1330_),
    .X(_0087_));
 sky130_fd_sc_hd__a21oi_1 _4890_ (.A1(_0420_),
    .A2(_0428_),
    .B1(_0412_),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_0412_),
    .B(_0637_),
    .Y(_1372_));
 sky130_fd_sc_hd__nor2_1 _4892_ (.A(_0430_),
    .B(_1371_),
    .Y(_1373_));
 sky130_fd_sc_hd__nor2_1 _4893_ (.A(_0646_),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__a32o_1 _4894_ (.A1(_0638_),
    .A2(_0646_),
    .A3(_1372_),
    .B1(_0570_),
    .B2(_0528_),
    .X(_1375_));
 sky130_fd_sc_hd__o221a_1 _4895_ (.A1(net132),
    .A2(_0622_),
    .B1(_1374_),
    .B2(_1375_),
    .C1(_0625_),
    .X(_1376_));
 sky130_fd_sc_hd__nor2_1 _4896_ (.A(_0625_),
    .B(_1373_),
    .Y(_1377_));
 sky130_fd_sc_hd__or3_4 _4897_ (.A(net83),
    .B(_1376_),
    .C(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__o21ai_1 _4898_ (.A1(\as1802.regs[2][0] ),
    .A2(net884),
    .B1(net851),
    .Y(_1379_));
 sky130_fd_sc_hd__a21o_1 _4899_ (.A1(_0706_),
    .A2(net885),
    .B1(net84),
    .X(_1380_));
 sky130_fd_sc_hd__xnor2_1 _4900_ (.A(_0739_),
    .B(_1355_),
    .Y(_1381_));
 sky130_fd_sc_hd__mux2_1 _4901_ (.A0(_0738_),
    .A1(_1381_),
    .S(net166),
    .X(_1382_));
 sky130_fd_sc_hd__nor2_1 _4902_ (.A(_0730_),
    .B(_0739_),
    .Y(_1383_));
 sky130_fd_sc_hd__o32a_1 _4903_ (.A1(_0740_),
    .A2(_0806_),
    .A3(_1383_),
    .B1(_1382_),
    .B2(_0573_),
    .X(_1384_));
 sky130_fd_sc_hd__o21a_1 _4904_ (.A1(_1358_),
    .A2(_1381_),
    .B1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(net154),
    .B(_0664_),
    .Y(_1386_));
 sky130_fd_sc_hd__o211a_1 _4906_ (.A1(_0661_),
    .A2(_1385_),
    .B1(_1386_),
    .C1(_0658_),
    .X(_1387_));
 sky130_fd_sc_hd__a211o_1 _4907_ (.A1(net82),
    .A2(_1382_),
    .B1(_1387_),
    .C1(_0676_),
    .X(_1388_));
 sky130_fd_sc_hd__nand2_1 _4908_ (.A(net23),
    .B(_0676_),
    .Y(_1389_));
 sky130_fd_sc_hd__o21ai_1 _4909_ (.A1(_0872_),
    .A2(_0891_),
    .B1(_0821_),
    .Y(_1390_));
 sky130_fd_sc_hd__o221a_1 _4910_ (.A1(_0412_),
    .A2(_0821_),
    .B1(_0892_),
    .B2(_1390_),
    .C1(net81),
    .X(_1391_));
 sky130_fd_sc_hd__a31o_1 _4911_ (.A1(net80),
    .A2(_1388_),
    .A3(_1389_),
    .B1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__o21ai_4 _4912_ (.A1(_0687_),
    .A2(_1392_),
    .B1(_1380_),
    .Y(_1393_));
 sky130_fd_sc_hd__mux2_1 _4913_ (.A0(net549),
    .A1(_1393_),
    .S(_1334_),
    .X(_1394_));
 sky130_fd_sc_hd__mux2_1 _4914_ (.A0(_1394_),
    .A1(_1378_),
    .S(_1330_),
    .X(_0088_));
 sky130_fd_sc_hd__nor2_1 _4915_ (.A(_0404_),
    .B(_0430_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_0404_),
    .B(_0638_),
    .Y(_1396_));
 sky130_fd_sc_hd__and2_1 _4917_ (.A(_0639_),
    .B(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_1 _4918_ (.A(_0622_),
    .B(_0646_),
    .Y(_1398_));
 sky130_fd_sc_hd__o22a_1 _4919_ (.A1(net130),
    .A2(_0622_),
    .B1(_1397_),
    .B2(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__o32a_1 _4920_ (.A1(_0431_),
    .A2(_0647_),
    .A3(_1395_),
    .B1(_1399_),
    .B2(_0624_),
    .X(_1400_));
 sky130_fd_sc_hd__or2_4 _4921_ (.A(net83),
    .B(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__nand2_1 _4922_ (.A(_0750_),
    .B(_0800_),
    .Y(_1402_));
 sky130_fd_sc_hd__a21oi_1 _4923_ (.A1(_0739_),
    .A2(_1355_),
    .B1(_0749_),
    .Y(_1403_));
 sky130_fd_sc_hd__a21o_1 _4924_ (.A1(_0750_),
    .A2(_0800_),
    .B1(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__o21a_1 _4925_ (.A1(_0729_),
    .A2(_0738_),
    .B1(_0748_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(_0748_),
    .A1(_1404_),
    .S(net166),
    .X(_1406_));
 sky130_fd_sc_hd__o32a_1 _4927_ (.A1(_0750_),
    .A2(_0806_),
    .A3(_1405_),
    .B1(_1406_),
    .B2(_0573_),
    .X(_1407_));
 sky130_fd_sc_hd__o21a_1 _4928_ (.A1(_1358_),
    .A2(_1404_),
    .B1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__o2bb2a_1 _4929_ (.A1_N(net151),
    .A2_N(_0664_),
    .B1(_1408_),
    .B2(_0661_),
    .X(_1409_));
 sky130_fd_sc_hd__mux2_1 _4930_ (.A0(_1406_),
    .A1(_1409_),
    .S(_0658_),
    .X(_1410_));
 sky130_fd_sc_hd__nor2_1 _4931_ (.A(net24),
    .B(net78),
    .Y(_1411_));
 sky130_fd_sc_hd__a211o_1 _4932_ (.A1(net78),
    .A2(_1410_),
    .B1(_1411_),
    .C1(net81),
    .X(_1412_));
 sky130_fd_sc_hd__xnor2_1 _4933_ (.A(_0893_),
    .B(_0894_),
    .Y(_1413_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(_0404_),
    .A1(_1413_),
    .S(_0821_),
    .X(_1414_));
 sky130_fd_sc_hd__o211a_1 _4935_ (.A1(net80),
    .A2(_1414_),
    .B1(_1412_),
    .C1(net84),
    .X(_1415_));
 sky130_fd_sc_hd__a21oi_2 _4936_ (.A1(\as1802.regs[2][3] ),
    .A2(_0706_),
    .B1(net84),
    .Y(_1416_));
 sky130_fd_sc_hd__a21oi_4 _4937_ (.A1(_0707_),
    .A2(_1416_),
    .B1(_1415_),
    .Y(_1417_));
 sky130_fd_sc_hd__mux2_1 _4938_ (.A0(net794),
    .A1(_1417_),
    .S(_1334_),
    .X(_1418_));
 sky130_fd_sc_hd__mux2_1 _4939_ (.A0(_1418_),
    .A1(_1401_),
    .S(_1330_),
    .X(_0089_));
 sky130_fd_sc_hd__nor2_1 _4940_ (.A(_0396_),
    .B(_0431_),
    .Y(_1419_));
 sky130_fd_sc_hd__nor2_1 _4941_ (.A(_0432_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(_0640_),
    .B(_0646_),
    .Y(_1421_));
 sky130_fd_sc_hd__a21o_1 _4943_ (.A1(_0396_),
    .A2(_0639_),
    .B1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__o211ai_1 _4944_ (.A1(_0646_),
    .A2(_1420_),
    .B1(_1422_),
    .C1(_0622_),
    .Y(_1423_));
 sky130_fd_sc_hd__or2_1 _4945_ (.A(net127),
    .B(_0622_),
    .X(_1424_));
 sky130_fd_sc_hd__nor2_1 _4946_ (.A(_0625_),
    .B(_1420_),
    .Y(_1425_));
 sky130_fd_sc_hd__a311o_4 _4947_ (.A1(_0625_),
    .A2(_1423_),
    .A3(_1424_),
    .B1(_1425_),
    .C1(net83),
    .X(_1426_));
 sky130_fd_sc_hd__xnor2_1 _4948_ (.A(net873),
    .B(_0707_),
    .Y(_1427_));
 sky130_fd_sc_hd__or2_1 _4949_ (.A(_0760_),
    .B(_0799_),
    .X(_1428_));
 sky130_fd_sc_hd__a21bo_1 _4950_ (.A1(_0758_),
    .A2(_1402_),
    .B1_N(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__inv_2 _4951_ (.A(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__a21o_1 _4952_ (.A1(net148),
    .A2(_0661_),
    .B1(net82),
    .X(_1431_));
 sky130_fd_sc_hd__nand2_1 _4953_ (.A(_0572_),
    .B(_1335_),
    .Y(_1432_));
 sky130_fd_sc_hd__o221a_1 _4954_ (.A1(net148),
    .A2(_0663_),
    .B1(_0759_),
    .B2(_1432_),
    .C1(_0662_),
    .X(_1433_));
 sky130_fd_sc_hd__xnor2_1 _4955_ (.A(_0750_),
    .B(_0758_),
    .Y(_1434_));
 sky130_fd_sc_hd__mux2_1 _4956_ (.A0(_0758_),
    .A1(_1429_),
    .S(net166),
    .X(_1435_));
 sky130_fd_sc_hd__o21a_1 _4957_ (.A1(_0573_),
    .A2(_1335_),
    .B1(_0806_),
    .X(_1436_));
 sky130_fd_sc_hd__o221a_1 _4958_ (.A1(_1358_),
    .A2(_1430_),
    .B1(_1434_),
    .B2(_1436_),
    .C1(_1433_),
    .X(_1437_));
 sky130_fd_sc_hd__o2bb2a_1 _4959_ (.A1_N(net82),
    .A2_N(_1435_),
    .B1(_1437_),
    .B2(_1431_),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_1 _4960_ (.A0(net25),
    .A1(_1438_),
    .S(net78),
    .X(_1439_));
 sky130_fd_sc_hd__a21oi_1 _4961_ (.A1(_0852_),
    .A2(_0895_),
    .B1(_0820_),
    .Y(_1440_));
 sky130_fd_sc_hd__a2bb2o_1 _4962_ (.A1_N(_0396_),
    .A2_N(_0821_),
    .B1(_0896_),
    .B2(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _4963_ (.A0(_1439_),
    .A1(_1441_),
    .S(net81),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_8 _4964_ (.A0(_1427_),
    .A1(_1442_),
    .S(net84),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _4965_ (.A0(net387),
    .A1(_1443_),
    .S(_1334_),
    .X(_1444_));
 sky130_fd_sc_hd__mux2_1 _4966_ (.A0(net388),
    .A1(_1426_),
    .S(_1330_),
    .X(_0090_));
 sky130_fd_sc_hd__o21a_1 _4967_ (.A1(_0432_),
    .A2(_0646_),
    .B1(_1421_),
    .X(_1445_));
 sky130_fd_sc_hd__and2_1 _4968_ (.A(_0388_),
    .B(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__o21ai_1 _4969_ (.A1(_0388_),
    .A2(_1445_),
    .B1(_0622_),
    .Y(_1447_));
 sky130_fd_sc_hd__o221a_1 _4970_ (.A1(net126),
    .A2(_0622_),
    .B1(_1446_),
    .B2(_1447_),
    .C1(_0625_),
    .X(_1448_));
 sky130_fd_sc_hd__nor2_1 _4971_ (.A(_0388_),
    .B(_0432_),
    .Y(_1449_));
 sky130_fd_sc_hd__or2_1 _4972_ (.A(_0433_),
    .B(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__a211o_4 _4973_ (.A1(_0624_),
    .A2(_1450_),
    .B1(_1448_),
    .C1(net83),
    .X(_1451_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_0770_),
    .B(_0800_),
    .Y(_1452_));
 sky130_fd_sc_hd__a22o_1 _4975_ (.A1(_0770_),
    .A2(_0800_),
    .B1(_1428_),
    .B2(_0768_),
    .X(_1453_));
 sky130_fd_sc_hd__or4_1 _4976_ (.A(net82),
    .B(_0661_),
    .C(_1358_),
    .D(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__and2_1 _4977_ (.A(_0760_),
    .B(_0768_),
    .X(_1455_));
 sky130_fd_sc_hd__o32a_1 _4978_ (.A1(_0770_),
    .A2(_1436_),
    .A3(_1455_),
    .B1(_1432_),
    .B2(_0768_),
    .X(_1456_));
 sky130_fd_sc_hd__a21bo_1 _4979_ (.A1(net238),
    .A2(_0664_),
    .B1_N(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(net165),
    .B(_1453_),
    .Y(_1458_));
 sky130_fd_sc_hd__o211a_1 _4981_ (.A1(net165),
    .A2(_0769_),
    .B1(_1458_),
    .C1(net82),
    .X(_1459_));
 sky130_fd_sc_hd__or4b_1 _4982_ (.A(_0676_),
    .B(_1457_),
    .C(_1459_),
    .D_N(_1454_),
    .X(_1460_));
 sky130_fd_sc_hd__o21a_1 _4983_ (.A1(net26),
    .A2(net78),
    .B1(net80),
    .X(_1461_));
 sky130_fd_sc_hd__and2b_1 _4984_ (.A_N(_0851_),
    .B(_0896_),
    .X(_1462_));
 sky130_fd_sc_hd__xnor2_1 _4985_ (.A(_0841_),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2_1 _4986_ (.A0(_0388_),
    .A1(_1463_),
    .S(_0821_),
    .X(_1464_));
 sky130_fd_sc_hd__o2bb2a_1 _4987_ (.A1_N(_1460_),
    .A2_N(_1461_),
    .B1(_1464_),
    .B2(net80),
    .X(_1465_));
 sky130_fd_sc_hd__o21ai_1 _4988_ (.A1(\as1802.regs[2][4] ),
    .A2(_0707_),
    .B1(\as1802.regs[2][5] ),
    .Y(_1466_));
 sky130_fd_sc_hd__and3_1 _4989_ (.A(_0687_),
    .B(_0708_),
    .C(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__a21oi_4 _4990_ (.A1(net84),
    .A2(_1465_),
    .B1(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__mux2_1 _4991_ (.A0(net771),
    .A1(_1468_),
    .S(_1334_),
    .X(_1469_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(_1469_),
    .A1(_1451_),
    .S(_1330_),
    .X(_0091_));
 sky130_fd_sc_hd__xnor2_1 _4993_ (.A(_0441_),
    .B(_0641_),
    .Y(_1470_));
 sky130_fd_sc_hd__o221a_1 _4994_ (.A1(net123),
    .A2(_0622_),
    .B1(_0646_),
    .B2(_0492_),
    .C1(_0625_),
    .X(_1471_));
 sky130_fd_sc_hd__o21a_1 _4995_ (.A1(_1398_),
    .A2(_1470_),
    .B1(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__a211o_4 _4996_ (.A1(_0492_),
    .A2(_0624_),
    .B1(net83),
    .C1(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__nand2_1 _4997_ (.A(\as1802.regs[2][6] ),
    .B(_0708_),
    .Y(_1474_));
 sky130_fd_sc_hd__a21oi_1 _4998_ (.A1(_0709_),
    .A2(_1474_),
    .B1(net84),
    .Y(_1475_));
 sky130_fd_sc_hd__or2_1 _4999_ (.A(_0780_),
    .B(_0799_),
    .X(_1476_));
 sky130_fd_sc_hd__a21bo_1 _5000_ (.A1(_0778_),
    .A2(_1452_),
    .B1_N(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__or2_1 _5001_ (.A(_1358_),
    .B(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__or2_1 _5002_ (.A(_0770_),
    .B(_0779_),
    .X(_1479_));
 sky130_fd_sc_hd__nand2_1 _5003_ (.A(_0780_),
    .B(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__o22a_1 _5004_ (.A1(_0778_),
    .A2(_1432_),
    .B1(_1436_),
    .B2(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__a21oi_1 _5005_ (.A1(_1478_),
    .A2(_1481_),
    .B1(_0661_),
    .Y(_1482_));
 sky130_fd_sc_hd__a211o_1 _5006_ (.A1(net142),
    .A2(_0664_),
    .B1(_1482_),
    .C1(_0657_),
    .X(_1483_));
 sky130_fd_sc_hd__mux2_1 _5007_ (.A0(_0778_),
    .A1(_1477_),
    .S(net165),
    .X(_1484_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(net82),
    .B(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__a31o_1 _5009_ (.A1(net27),
    .A2(_0673_),
    .A3(_0675_),
    .B1(net81),
    .X(_1486_));
 sky130_fd_sc_hd__a31o_1 _5010_ (.A1(net78),
    .A2(_1483_),
    .A3(_1485_),
    .B1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__and2_1 _5011_ (.A(_0897_),
    .B(_0920_),
    .X(_1488_));
 sky130_fd_sc_hd__or2_1 _5012_ (.A(_0908_),
    .B(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__a21oi_1 _5013_ (.A1(_0908_),
    .A2(_1488_),
    .B1(_0820_),
    .Y(_1490_));
 sky130_fd_sc_hd__a221o_1 _5014_ (.A1(_0442_),
    .A2(_0820_),
    .B1(_1489_),
    .B2(_1490_),
    .C1(net80),
    .X(_1491_));
 sky130_fd_sc_hd__a31o_4 _5015_ (.A1(net84),
    .A2(_1487_),
    .A3(_1491_),
    .B1(_1475_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _5016_ (.A0(net641),
    .A1(_1492_),
    .S(_1334_),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _5017_ (.A0(net642),
    .A1(_1473_),
    .S(_1330_),
    .X(_0092_));
 sky130_fd_sc_hd__and2_1 _5018_ (.A(_0451_),
    .B(_0642_),
    .X(_1494_));
 sky130_fd_sc_hd__nor2_1 _5019_ (.A(_0643_),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__o22a_1 _5020_ (.A1(net120),
    .A2(_0622_),
    .B1(_1398_),
    .B2(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__o22a_1 _5021_ (.A1(_0490_),
    .A2(_0647_),
    .B1(_1496_),
    .B2(_0624_),
    .X(_1497_));
 sky130_fd_sc_hd__or2_4 _5022_ (.A(net83),
    .B(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__a21o_1 _5023_ (.A1(_0788_),
    .A2(_1476_),
    .B1(_0802_),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _5024_ (.A0(_0788_),
    .A1(_1499_),
    .S(net165),
    .X(_1500_));
 sky130_fd_sc_hd__o221a_1 _5025_ (.A1(_3478_),
    .A2(_0663_),
    .B1(_0788_),
    .B2(_1432_),
    .C1(_0662_),
    .X(_1501_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_0780_),
    .B(_0788_),
    .Y(_1502_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_0790_),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__o221a_1 _5028_ (.A1(_1358_),
    .A2(_1499_),
    .B1(_1503_),
    .B2(_1436_),
    .C1(_1501_),
    .X(_1504_));
 sky130_fd_sc_hd__a211o_1 _5029_ (.A1(_3478_),
    .A2(_0661_),
    .B1(_1504_),
    .C1(net82),
    .X(_1505_));
 sky130_fd_sc_hd__o21ai_1 _5030_ (.A1(_0658_),
    .A2(_1500_),
    .B1(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(net28),
    .A1(_1506_),
    .S(net78),
    .X(_1507_));
 sky130_fd_sc_hd__and3b_1 _5032_ (.A_N(_0917_),
    .B(_1489_),
    .C(_0907_),
    .X(_1508_));
 sky130_fd_sc_hd__a21boi_1 _5033_ (.A1(_0907_),
    .A2(_1489_),
    .B1_N(_0917_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_0451_),
    .B(_0820_),
    .Y(_1510_));
 sky130_fd_sc_hd__o311a_1 _5035_ (.A1(_0820_),
    .A2(_1508_),
    .A3(_1509_),
    .B1(_1510_),
    .C1(net81),
    .X(_1511_));
 sky130_fd_sc_hd__a211o_1 _5036_ (.A1(net80),
    .A2(_1507_),
    .B1(_1511_),
    .C1(_0687_),
    .X(_1512_));
 sky130_fd_sc_hd__and2_1 _5037_ (.A(net842),
    .B(_0709_),
    .X(_1513_));
 sky130_fd_sc_hd__o31a_4 _5038_ (.A1(net85),
    .A2(_0710_),
    .A3(_1513_),
    .B1(_1512_),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_1 _5039_ (.A0(net784),
    .A1(_1514_),
    .S(_1334_),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _5040_ (.A0(net785),
    .A1(_1498_),
    .S(_1330_),
    .X(_0093_));
 sky130_fd_sc_hd__and3_4 _5041_ (.A(_1271_),
    .B(_1294_),
    .C(_1329_),
    .X(_1516_));
 sky130_fd_sc_hd__and3_4 _5042_ (.A(_1274_),
    .B(_1296_),
    .C(_1333_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _5043_ (.A0(net538),
    .A1(_1347_),
    .S(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_1 _5044_ (.A0(net539),
    .A1(_1332_),
    .S(_1516_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _5045_ (.A0(net814),
    .A1(_1369_),
    .S(_1517_),
    .X(_1519_));
 sky130_fd_sc_hd__mux2_1 _5046_ (.A0(net815),
    .A1(_1353_),
    .S(_1516_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _5047_ (.A0(net768),
    .A1(_1393_),
    .S(_1517_),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_1 _5048_ (.A0(_1520_),
    .A1(_1378_),
    .S(_1516_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(net474),
    .A1(_1417_),
    .S(_1517_),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _5050_ (.A0(_1521_),
    .A1(_1401_),
    .S(_1516_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _5051_ (.A0(net527),
    .A1(_1443_),
    .S(_1517_),
    .X(_1522_));
 sky130_fd_sc_hd__mux2_1 _5052_ (.A0(net528),
    .A1(_1426_),
    .S(_1516_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _5053_ (.A0(net468),
    .A1(_1468_),
    .S(_1517_),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _5054_ (.A0(_1523_),
    .A1(_1451_),
    .S(_1516_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(net478),
    .A1(_1492_),
    .S(_1517_),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _5056_ (.A0(net479),
    .A1(_1473_),
    .S(_1516_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(net517),
    .A1(_1514_),
    .S(_1517_),
    .X(_1525_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(net518),
    .A1(_1498_),
    .S(_1516_),
    .X(_0101_));
 sky130_fd_sc_hd__and3b_4 _5059_ (.A_N(_0633_),
    .B(_1270_),
    .C(_1329_),
    .X(_1526_));
 sky130_fd_sc_hd__and3_4 _5060_ (.A(_0702_),
    .B(_1273_),
    .C(_1333_),
    .X(_1527_));
 sky130_fd_sc_hd__mux2_1 _5061_ (.A0(net773),
    .A1(_1347_),
    .S(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _5062_ (.A0(net774),
    .A1(_1332_),
    .S(_1526_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _5063_ (.A0(net595),
    .A1(_1369_),
    .S(_1527_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _5064_ (.A0(net596),
    .A1(_1353_),
    .S(_1526_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _5065_ (.A0(net630),
    .A1(_1393_),
    .S(_1527_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(_1530_),
    .A1(_1378_),
    .S(_1526_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(net829),
    .A1(_1417_),
    .S(_1527_),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _5068_ (.A0(_1531_),
    .A1(_1401_),
    .S(_1526_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(net470),
    .A1(_1443_),
    .S(_1527_),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(net471),
    .A1(_1426_),
    .S(_1526_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _5071_ (.A0(net782),
    .A1(_1468_),
    .S(_1527_),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_1 _5072_ (.A0(_1533_),
    .A1(_1451_),
    .S(_1526_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _5073_ (.A0(net497),
    .A1(_1492_),
    .S(_1527_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_1 _5074_ (.A0(_1534_),
    .A1(_1473_),
    .S(_1526_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _5075_ (.A0(net394),
    .A1(_1514_),
    .S(_1527_),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(net395),
    .A1(_1498_),
    .S(_1526_),
    .X(_0109_));
 sky130_fd_sc_hd__and3_4 _5077_ (.A(_1294_),
    .B(_1316_),
    .C(_1329_),
    .X(_1536_));
 sky130_fd_sc_hd__and3_4 _5078_ (.A(_1296_),
    .B(_1318_),
    .C(_1333_),
    .X(_1537_));
 sky130_fd_sc_hd__mux2_1 _5079_ (.A0(net577),
    .A1(_1347_),
    .S(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__mux2_1 _5080_ (.A0(net578),
    .A1(_1332_),
    .S(_1536_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _5081_ (.A0(net798),
    .A1(_1369_),
    .S(_1537_),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_1 _5082_ (.A0(net799),
    .A1(_1353_),
    .S(_1536_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _5083_ (.A0(net775),
    .A1(_1393_),
    .S(_1537_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _5084_ (.A0(_1540_),
    .A1(_1378_),
    .S(_1536_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5085_ (.A0(net516),
    .A1(_1417_),
    .S(_1537_),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _5086_ (.A0(_1541_),
    .A1(_1401_),
    .S(_1536_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5087_ (.A0(net550),
    .A1(_1443_),
    .S(_1537_),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _5088_ (.A0(net551),
    .A1(_1426_),
    .S(_1536_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _5089_ (.A0(net381),
    .A1(_1468_),
    .S(_1537_),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _5090_ (.A0(_1543_),
    .A1(_1451_),
    .S(_1536_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(net402),
    .A1(_1492_),
    .S(_1537_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _5092_ (.A0(net403),
    .A1(_1473_),
    .S(_1536_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(net416),
    .A1(_1514_),
    .S(_1537_),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _5094_ (.A0(net417),
    .A1(_1498_),
    .S(_1536_),
    .X(_0117_));
 sky130_fd_sc_hd__and3_4 _5095_ (.A(_1257_),
    .B(_1270_),
    .C(_1329_),
    .X(_1546_));
 sky130_fd_sc_hd__and3_4 _5096_ (.A(_1260_),
    .B(_1273_),
    .C(_1333_),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(net839),
    .A1(_1347_),
    .S(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _5098_ (.A0(_1548_),
    .A1(_1332_),
    .S(_1546_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _5099_ (.A0(net836),
    .A1(_1369_),
    .S(_1547_),
    .X(_1549_));
 sky130_fd_sc_hd__mux2_1 _5100_ (.A0(net837),
    .A1(_1353_),
    .S(_1546_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5101_ (.A0(net851),
    .A1(_1393_),
    .S(_1547_),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_1 _5102_ (.A0(_1550_),
    .A1(_1378_),
    .S(_1546_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5103_ (.A0(net857),
    .A1(_1417_),
    .S(_1547_),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_1 _5104_ (.A0(_1551_),
    .A1(_1401_),
    .S(_1546_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(net873),
    .A1(_1443_),
    .S(_1547_),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(_1552_),
    .A1(_1426_),
    .S(_1546_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(net847),
    .A1(_1468_),
    .S(_1547_),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(_1553_),
    .A1(_1451_),
    .S(_1546_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _5109_ (.A0(net841),
    .A1(_1492_),
    .S(_1547_),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(_1554_),
    .A1(_1473_),
    .S(_1546_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(net842),
    .A1(_1514_),
    .S(_1547_),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _5112_ (.A0(_1555_),
    .A1(_1498_),
    .S(_1546_),
    .X(_0125_));
 sky130_fd_sc_hd__and3_4 _5113_ (.A(_1270_),
    .B(_1316_),
    .C(_1329_),
    .X(_1556_));
 sky130_fd_sc_hd__and3_4 _5114_ (.A(_1273_),
    .B(_1318_),
    .C(_1333_),
    .X(_1557_));
 sky130_fd_sc_hd__mux2_1 _5115_ (.A0(net606),
    .A1(_1347_),
    .S(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _5116_ (.A0(net607),
    .A1(_1332_),
    .S(_1556_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(net495),
    .A1(_1369_),
    .S(_1557_),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(net496),
    .A1(_1353_),
    .S(_1556_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5119_ (.A0(net591),
    .A1(_1393_),
    .S(_1557_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _5120_ (.A0(_1560_),
    .A1(_1378_),
    .S(_1556_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5121_ (.A0(net801),
    .A1(_1417_),
    .S(_1557_),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _5122_ (.A0(_1561_),
    .A1(_1401_),
    .S(_1556_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(net428),
    .A1(_1443_),
    .S(_1557_),
    .X(_1562_));
 sky130_fd_sc_hd__mux2_1 _5124_ (.A0(_1562_),
    .A1(_1426_),
    .S(_1556_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _5125_ (.A0(net759),
    .A1(_1468_),
    .S(_1557_),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_1 _5126_ (.A0(_1563_),
    .A1(_1451_),
    .S(_1556_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(net583),
    .A1(_1492_),
    .S(_1557_),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_1 _5128_ (.A0(_1564_),
    .A1(_1473_),
    .S(_1556_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(net786),
    .A1(_1514_),
    .S(_1557_),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_1 _5130_ (.A0(net787),
    .A1(_1498_),
    .S(_1556_),
    .X(_0133_));
 sky130_fd_sc_hd__nor3_2 _5131_ (.A(_3463_),
    .B(net366),
    .C(_3544_),
    .Y(_1566_));
 sky130_fd_sc_hd__or3_4 _5132_ (.A(_3463_),
    .B(net366),
    .C(_3544_),
    .X(_1567_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_3444_),
    .B(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__o211a_1 _5134_ (.A1(net31),
    .A2(_1567_),
    .B1(_1568_),
    .C1(net207),
    .X(_0134_));
 sky130_fd_sc_hd__or2_1 _5135_ (.A(net169),
    .B(_1566_),
    .X(_1569_));
 sky130_fd_sc_hd__o211a_1 _5136_ (.A1(net32),
    .A2(_1567_),
    .B1(_1569_),
    .C1(net207),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _5137_ (.A0(net167),
    .A1(net33),
    .S(_1566_),
    .X(_1570_));
 sky130_fd_sc_hd__or2_1 _5138_ (.A(net206),
    .B(_1570_),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_1 _5139_ (.A(net117),
    .B(_1567_),
    .Y(_1571_));
 sky130_fd_sc_hd__o211a_1 _5140_ (.A1(net34),
    .A2(_1567_),
    .B1(_1571_),
    .C1(net207),
    .X(_0137_));
 sky130_fd_sc_hd__or3b_4 _5141_ (.A(_0630_),
    .B(_1328_),
    .C_N(_1257_),
    .X(_1572_));
 sky130_fd_sc_hd__and3_4 _5142_ (.A(_0694_),
    .B(_1260_),
    .C(_1333_),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _5143_ (.A0(net698),
    .A1(_1347_),
    .S(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _5144_ (.A0(_1332_),
    .A1(net699),
    .S(_1572_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _5145_ (.A0(net682),
    .A1(_1369_),
    .S(_1573_),
    .X(_1575_));
 sky130_fd_sc_hd__mux2_1 _5146_ (.A0(_1353_),
    .A1(net683),
    .S(_1572_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(net720),
    .A1(_1393_),
    .S(_1573_),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_1 _5148_ (.A0(_1378_),
    .A1(net721),
    .S(_1572_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _5149_ (.A0(net816),
    .A1(_1417_),
    .S(_1573_),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_1 _5150_ (.A0(_1401_),
    .A1(_1577_),
    .S(_1572_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(net778),
    .A1(_1443_),
    .S(_1573_),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _5152_ (.A0(_1426_),
    .A1(net779),
    .S(_1572_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(net564),
    .A1(_1468_),
    .S(_1573_),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_1 _5154_ (.A0(_1451_),
    .A1(_1579_),
    .S(_1572_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(net803),
    .A1(_1492_),
    .S(_1573_),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _5156_ (.A0(_1473_),
    .A1(net804),
    .S(_1572_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(net765),
    .A1(_1514_),
    .S(_1573_),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_1 _5158_ (.A0(_1498_),
    .A1(net766),
    .S(_1572_),
    .X(_0145_));
 sky130_fd_sc_hd__and3_4 _5159_ (.A(_0635_),
    .B(_1271_),
    .C(_1294_),
    .X(_1582_));
 sky130_fd_sc_hd__and3_4 _5160_ (.A(_0704_),
    .B(_1274_),
    .C(_1296_),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(net409),
    .A1(_0926_),
    .S(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__mux2_1 _5162_ (.A0(net410),
    .A1(_0652_),
    .S(_1582_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _5163_ (.A0(net489),
    .A1(_0974_),
    .S(_1583_),
    .X(_1585_));
 sky130_fd_sc_hd__mux2_1 _5164_ (.A0(_1585_),
    .A1(_0934_),
    .S(_1582_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(net707),
    .A1(_1022_),
    .S(_1583_),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _5166_ (.A0(net708),
    .A1(_0982_),
    .S(_1582_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _5167_ (.A0(net440),
    .A1(_1067_),
    .S(_1583_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(net441),
    .A1(_1030_),
    .S(_1582_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _5169_ (.A0(net543),
    .A1(_1117_),
    .S(_1583_),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_1 _5170_ (.A0(_1588_),
    .A1(_1075_),
    .S(_1582_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _5171_ (.A0(net694),
    .A1(_1165_),
    .S(_1583_),
    .X(_1589_));
 sky130_fd_sc_hd__mux2_1 _5172_ (.A0(net695),
    .A1(_1125_),
    .S(_1582_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5173_ (.A0(net447),
    .A1(_1214_),
    .S(_1583_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _5174_ (.A0(_1590_),
    .A1(_1172_),
    .S(_1582_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5175_ (.A0(net540),
    .A1(_1253_),
    .S(_1583_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _5176_ (.A0(_1591_),
    .A1(_1219_),
    .S(_1582_),
    .X(_0153_));
 sky130_fd_sc_hd__or3_4 _5177_ (.A(_0630_),
    .B(_0633_),
    .C(_1328_),
    .X(_1592_));
 sky130_fd_sc_hd__and3_4 _5178_ (.A(_0694_),
    .B(_0702_),
    .C(_1333_),
    .X(_1593_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(net749),
    .A1(_1347_),
    .S(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _5180_ (.A0(_1332_),
    .A1(net750),
    .S(_1592_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(net780),
    .A1(_1369_),
    .S(_1593_),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_1 _5182_ (.A0(_1353_),
    .A1(net781),
    .S(_1592_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5183_ (.A0(net574),
    .A1(_1393_),
    .S(_1593_),
    .X(_1596_));
 sky130_fd_sc_hd__mux2_1 _5184_ (.A0(_1378_),
    .A1(net575),
    .S(_1592_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _5185_ (.A0(net627),
    .A1(_1417_),
    .S(_1593_),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _5186_ (.A0(_1401_),
    .A1(_1597_),
    .S(_1592_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _5187_ (.A0(net661),
    .A1(_1443_),
    .S(_1593_),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_1 _5188_ (.A0(_1426_),
    .A1(net662),
    .S(_1592_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(net738),
    .A1(_1468_),
    .S(_1593_),
    .X(_1599_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(_1451_),
    .A1(_1599_),
    .S(_1592_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(net544),
    .A1(_1492_),
    .S(_1593_),
    .X(_1600_));
 sky130_fd_sc_hd__mux2_1 _5192_ (.A0(_1473_),
    .A1(net545),
    .S(_1592_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(net510),
    .A1(_1514_),
    .S(_1593_),
    .X(_1601_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(_1498_),
    .A1(net511),
    .S(_1592_),
    .X(_0161_));
 sky130_fd_sc_hd__or3b_4 _5195_ (.A(_0630_),
    .B(_1328_),
    .C_N(_1316_),
    .X(_1602_));
 sky130_fd_sc_hd__and3_4 _5196_ (.A(_0694_),
    .B(_1318_),
    .C(_1333_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _5197_ (.A0(net744),
    .A1(_1347_),
    .S(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__mux2_1 _5198_ (.A0(_1332_),
    .A1(net745),
    .S(_1602_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(net755),
    .A1(_1369_),
    .S(_1603_),
    .X(_1605_));
 sky130_fd_sc_hd__mux2_1 _5200_ (.A0(_1353_),
    .A1(net756),
    .S(_1602_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(net475),
    .A1(_1393_),
    .S(_1603_),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(_1378_),
    .A1(net476),
    .S(_1602_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _5203_ (.A0(net620),
    .A1(_1417_),
    .S(_1603_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _5204_ (.A0(_1401_),
    .A1(_1607_),
    .S(_1602_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5205_ (.A0(net579),
    .A1(_1443_),
    .S(_1603_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_1 _5206_ (.A0(_1426_),
    .A1(net580),
    .S(_1602_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5207_ (.A0(net633),
    .A1(_1468_),
    .S(_1603_),
    .X(_1609_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(_1451_),
    .A1(_1609_),
    .S(_1602_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5209_ (.A0(net806),
    .A1(_1492_),
    .S(_1603_),
    .X(_1610_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(_1473_),
    .A1(net807),
    .S(_1602_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(net541),
    .A1(_1514_),
    .S(_1603_),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(_1498_),
    .A1(net542),
    .S(_1602_),
    .X(_0169_));
 sky130_fd_sc_hd__and3b_4 _5213_ (.A_N(_0630_),
    .B(_1271_),
    .C(_1329_),
    .X(_1612_));
 sky130_fd_sc_hd__and3_4 _5214_ (.A(_0694_),
    .B(_1274_),
    .C(_1333_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _5215_ (.A0(net615),
    .A1(_1347_),
    .S(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(net616),
    .A1(_1332_),
    .S(_1612_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5217_ (.A0(net696),
    .A1(_1369_),
    .S(_1613_),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_1 _5218_ (.A0(net697),
    .A1(_1353_),
    .S(_1612_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(net586),
    .A1(_1393_),
    .S(_1613_),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_1 _5220_ (.A0(net587),
    .A1(_1378_),
    .S(_1612_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(net735),
    .A1(_1417_),
    .S(_1613_),
    .X(_1617_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(_1617_),
    .A1(_1401_),
    .S(_1612_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5223_ (.A0(net700),
    .A1(_1443_),
    .S(_1613_),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_1 _5224_ (.A0(net701),
    .A1(_1426_),
    .S(_1612_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5225_ (.A0(net599),
    .A1(_1468_),
    .S(_1613_),
    .X(_1619_));
 sky130_fd_sc_hd__mux2_1 _5226_ (.A0(_1619_),
    .A1(_1451_),
    .S(_1612_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5227_ (.A0(net601),
    .A1(_1492_),
    .S(_1613_),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _5228_ (.A0(net602),
    .A1(_1473_),
    .S(_1612_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5229_ (.A0(net592),
    .A1(_1514_),
    .S(_1613_),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_1 _5230_ (.A0(net593),
    .A1(_1498_),
    .S(_1612_),
    .X(_0177_));
 sky130_fd_sc_hd__or3b_4 _5231_ (.A(_0633_),
    .B(_1328_),
    .C_N(_1256_),
    .X(_1622_));
 sky130_fd_sc_hd__and3_4 _5232_ (.A(_0702_),
    .B(_1259_),
    .C(_1333_),
    .X(_1623_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(net761),
    .A1(_1347_),
    .S(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _5234_ (.A0(_1332_),
    .A1(net762),
    .S(_1622_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(net757),
    .A1(_1369_),
    .S(_1623_),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_1 _5236_ (.A0(_1353_),
    .A1(net758),
    .S(_1622_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _5237_ (.A0(net492),
    .A1(_1393_),
    .S(_1623_),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_1 _5238_ (.A0(_1378_),
    .A1(net493),
    .S(_1622_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _5239_ (.A0(net802),
    .A1(_1417_),
    .S(_1623_),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(_1401_),
    .A1(_1627_),
    .S(_1622_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(net730),
    .A1(_1443_),
    .S(_1623_),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(_1426_),
    .A1(net731),
    .S(_1622_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(net716),
    .A1(_1468_),
    .S(_1623_),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(_1451_),
    .A1(_1629_),
    .S(_1622_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _5245_ (.A0(net723),
    .A1(_1492_),
    .S(_1623_),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _5246_ (.A0(_1473_),
    .A1(net724),
    .S(_1622_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(net753),
    .A1(_1514_),
    .S(_1623_),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(_1498_),
    .A1(net754),
    .S(_1622_),
    .X(_0185_));
 sky130_fd_sc_hd__and3_4 _5249_ (.A(_1256_),
    .B(_1257_),
    .C(_1329_),
    .X(_1632_));
 sky130_fd_sc_hd__and3_4 _5250_ (.A(_1259_),
    .B(_1260_),
    .C(_1333_),
    .X(_1633_));
 sky130_fd_sc_hd__mux2_1 _5251_ (.A0(net452),
    .A1(_1347_),
    .S(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(net453),
    .A1(_1332_),
    .S(_1632_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _5253_ (.A0(net504),
    .A1(_1369_),
    .S(_1633_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(net505),
    .A1(_1353_),
    .S(_1632_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _5255_ (.A0(net552),
    .A1(_1393_),
    .S(_1633_),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(net553),
    .A1(_1378_),
    .S(_1632_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(net740),
    .A1(_1417_),
    .S(_1633_),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(_1637_),
    .A1(_1401_),
    .S(_1632_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _5259_ (.A0(net536),
    .A1(_1443_),
    .S(_1633_),
    .X(_1638_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(net537),
    .A1(_1426_),
    .S(_1632_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _5261_ (.A0(net608),
    .A1(_1468_),
    .S(_1633_),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(_1639_),
    .A1(_1451_),
    .S(_1632_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(net420),
    .A1(_1492_),
    .S(_1633_),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(_1640_),
    .A1(_1473_),
    .S(_1632_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5265_ (.A0(net506),
    .A1(_1514_),
    .S(_1633_),
    .X(_1641_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(net507),
    .A1(_1498_),
    .S(_1632_),
    .X(_0193_));
 sky130_fd_sc_hd__and3_4 _5267_ (.A(_1270_),
    .B(_1271_),
    .C(_1329_),
    .X(_1642_));
 sky130_fd_sc_hd__and3_4 _5268_ (.A(_1273_),
    .B(_1274_),
    .C(_1333_),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(net705),
    .A1(_1347_),
    .S(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__mux2_1 _5270_ (.A0(net706),
    .A1(_1332_),
    .S(_1642_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _5271_ (.A0(net612),
    .A1(_1369_),
    .S(_1643_),
    .X(_1645_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net613),
    .A1(_1353_),
    .S(_1642_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5273_ (.A0(net795),
    .A1(_1393_),
    .S(_1643_),
    .X(_1646_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(_1646_),
    .A1(_1378_),
    .S(_1642_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(net680),
    .A1(_1417_),
    .S(_1643_),
    .X(_1647_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(_1647_),
    .A1(_1401_),
    .S(_1642_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(net646),
    .A1(_1443_),
    .S(_1643_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(net647),
    .A1(_1426_),
    .S(_1642_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(net622),
    .A1(_1468_),
    .S(_1643_),
    .X(_1649_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(_1649_),
    .A1(_1451_),
    .S(_1642_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(net664),
    .A1(_1492_),
    .S(_1643_),
    .X(_1650_));
 sky130_fd_sc_hd__mux2_1 _5282_ (.A0(_1650_),
    .A1(_1473_),
    .S(_1642_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(net709),
    .A1(_1514_),
    .S(_1643_),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(net710),
    .A1(_1498_),
    .S(_1642_),
    .X(_0201_));
 sky130_fd_sc_hd__and3_4 _5285_ (.A(_1256_),
    .B(_1316_),
    .C(_1329_),
    .X(_1652_));
 sky130_fd_sc_hd__and3_4 _5286_ (.A(_1259_),
    .B(_1318_),
    .C(_1333_),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(net426),
    .A1(_1347_),
    .S(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_1 _5288_ (.A0(net427),
    .A1(_1332_),
    .S(_1652_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(net512),
    .A1(_1369_),
    .S(_1653_),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(net513),
    .A1(_1353_),
    .S(_1652_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(net486),
    .A1(_1393_),
    .S(_1653_),
    .X(_1656_));
 sky130_fd_sc_hd__mux2_1 _5292_ (.A0(net487),
    .A1(_1378_),
    .S(_1652_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(net660),
    .A1(_1417_),
    .S(_1653_),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(_1657_),
    .A1(_1401_),
    .S(_1652_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(net702),
    .A1(_1443_),
    .S(_1653_),
    .X(_1658_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(net703),
    .A1(_1426_),
    .S(_1652_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(net502),
    .A1(_1468_),
    .S(_1653_),
    .X(_1659_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(_1659_),
    .A1(_1451_),
    .S(_1652_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(net414),
    .A1(_1492_),
    .S(_1653_),
    .X(_1660_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net415),
    .A1(_1473_),
    .S(_1652_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(net521),
    .A1(_1514_),
    .S(_1653_),
    .X(_1661_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(net522),
    .A1(_1498_),
    .S(_1652_),
    .X(_0209_));
 sky130_fd_sc_hd__and3_4 _5303_ (.A(_1256_),
    .B(_1271_),
    .C(_1329_),
    .X(_1662_));
 sky130_fd_sc_hd__and3_4 _5304_ (.A(_1259_),
    .B(_1274_),
    .C(_1333_),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(net617),
    .A1(_1347_),
    .S(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _5306_ (.A0(net618),
    .A1(_1332_),
    .S(_1662_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(net558),
    .A1(_1369_),
    .S(_1663_),
    .X(_1665_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net559),
    .A1(_1353_),
    .S(_1662_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net456),
    .A1(_1393_),
    .S(_1663_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net457),
    .A1(_1378_),
    .S(_1662_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(net555),
    .A1(_1417_),
    .S(_1663_),
    .X(_1667_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(_1667_),
    .A1(_1401_),
    .S(_1662_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5313_ (.A0(net747),
    .A1(_1443_),
    .S(_1663_),
    .X(_1668_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(net748),
    .A1(_1426_),
    .S(_1662_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(net637),
    .A1(_1468_),
    .S(_1663_),
    .X(_1669_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(_1669_),
    .A1(_1451_),
    .S(_1662_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5317_ (.A0(net450),
    .A1(_1492_),
    .S(_1663_),
    .X(_1670_));
 sky130_fd_sc_hd__mux2_1 _5318_ (.A0(net451),
    .A1(_1473_),
    .S(_1662_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(net404),
    .A1(_1514_),
    .S(_1663_),
    .X(_1671_));
 sky130_fd_sc_hd__mux2_1 _5320_ (.A0(net405),
    .A1(_1498_),
    .S(_1662_),
    .X(_0217_));
 sky130_fd_sc_hd__or3b_4 _5321_ (.A(_0633_),
    .B(_1328_),
    .C_N(_1294_),
    .X(_1672_));
 sky130_fd_sc_hd__and3_4 _5322_ (.A(_0702_),
    .B(_1296_),
    .C(_1333_),
    .X(_1673_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(net572),
    .A1(_1347_),
    .S(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(_1332_),
    .A1(net573),
    .S(_1672_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(net812),
    .A1(_1369_),
    .S(_1673_),
    .X(_1675_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(_1353_),
    .A1(net813),
    .S(_1672_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5327_ (.A0(net669),
    .A1(_1393_),
    .S(_1673_),
    .X(_1676_));
 sky130_fd_sc_hd__mux2_1 _5328_ (.A0(_1378_),
    .A1(_1676_),
    .S(_1672_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5329_ (.A0(net823),
    .A1(_1417_),
    .S(_1673_),
    .X(_1677_));
 sky130_fd_sc_hd__mux2_1 _5330_ (.A0(_1401_),
    .A1(_1677_),
    .S(_1672_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(net500),
    .A1(_1443_),
    .S(_1673_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(_1426_),
    .A1(net501),
    .S(_1672_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5333_ (.A0(net635),
    .A1(_1468_),
    .S(_1673_),
    .X(_1679_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(_1451_),
    .A1(_1679_),
    .S(_1672_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(net648),
    .A1(_1492_),
    .S(_1673_),
    .X(_1680_));
 sky130_fd_sc_hd__mux2_1 _5336_ (.A0(_1473_),
    .A1(net649),
    .S(_1672_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net769),
    .A1(_1514_),
    .S(_1673_),
    .X(_1681_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(_1498_),
    .A1(net770),
    .S(_1672_),
    .X(_0225_));
 sky130_fd_sc_hd__or3b_4 _5339_ (.A(_0630_),
    .B(_0634_),
    .C_N(_1257_),
    .X(_1682_));
 sky130_fd_sc_hd__and3_4 _5340_ (.A(_0694_),
    .B(_0704_),
    .C(_1260_),
    .X(_1683_));
 sky130_fd_sc_hd__mux2_1 _5341_ (.A0(net556),
    .A1(_0926_),
    .S(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(_0652_),
    .A1(net557),
    .S(_1682_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(net681),
    .A1(_0974_),
    .S(_1683_),
    .X(_1685_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(_0934_),
    .A1(_1685_),
    .S(_1682_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(net628),
    .A1(_1022_),
    .S(_1683_),
    .X(_1686_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(_0982_),
    .A1(net629),
    .S(_1682_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(net728),
    .A1(_1067_),
    .S(_1683_),
    .X(_1687_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(_1030_),
    .A1(net729),
    .S(_1682_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(net741),
    .A1(_1117_),
    .S(_1683_),
    .X(_1688_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(_1075_),
    .A1(_1688_),
    .S(_1682_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(net790),
    .A1(_1165_),
    .S(_1683_),
    .X(_1689_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(_1125_),
    .A1(net791),
    .S(_1682_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(net686),
    .A1(_1214_),
    .S(_1683_),
    .X(_1690_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(_1172_),
    .A1(_1690_),
    .S(_1682_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5355_ (.A0(net679),
    .A1(_1253_),
    .S(_1683_),
    .X(_1691_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(_1219_),
    .A1(_1691_),
    .S(_1682_),
    .X(_0233_));
 sky130_fd_sc_hd__or3b_4 _5357_ (.A(_0630_),
    .B(_0634_),
    .C_N(_1316_),
    .X(_1692_));
 sky130_fd_sc_hd__and3_4 _5358_ (.A(_0694_),
    .B(_0704_),
    .C(_1318_),
    .X(_1693_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(net763),
    .A1(_0926_),
    .S(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_1 _5360_ (.A0(_0652_),
    .A1(net764),
    .S(_1692_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net789),
    .A1(_0974_),
    .S(_1693_),
    .X(_1695_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(_0934_),
    .A1(_1695_),
    .S(_1692_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(net655),
    .A1(_1022_),
    .S(_1693_),
    .X(_1696_));
 sky130_fd_sc_hd__mux2_1 _5364_ (.A0(_0982_),
    .A1(net656),
    .S(_1692_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(net424),
    .A1(_1067_),
    .S(_1693_),
    .X(_1697_));
 sky130_fd_sc_hd__mux2_1 _5366_ (.A0(_1030_),
    .A1(net425),
    .S(_1692_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(net692),
    .A1(_1117_),
    .S(_1693_),
    .X(_1698_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(_1075_),
    .A1(_1698_),
    .S(_1692_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(net407),
    .A1(_1165_),
    .S(_1693_),
    .X(_1699_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(_1125_),
    .A1(net408),
    .S(_1692_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net523),
    .A1(_1214_),
    .S(_1693_),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(_1172_),
    .A1(_1700_),
    .S(_1692_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net519),
    .A1(_1253_),
    .S(_1693_),
    .X(_1701_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(_1219_),
    .A1(_1701_),
    .S(_1692_),
    .X(_0241_));
 sky130_fd_sc_hd__and3b_4 _5375_ (.A_N(_0630_),
    .B(_0635_),
    .C(_1271_),
    .X(_1702_));
 sky130_fd_sc_hd__and3_4 _5376_ (.A(_0694_),
    .B(_0704_),
    .C(_1274_),
    .X(_1703_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(net466),
    .A1(_0926_),
    .S(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__mux2_1 _5378_ (.A0(net467),
    .A1(_0652_),
    .S(_1702_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(net671),
    .A1(_0974_),
    .S(_1703_),
    .X(_1705_));
 sky130_fd_sc_hd__mux2_1 _5380_ (.A0(_1705_),
    .A1(_0934_),
    .S(_1702_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(net667),
    .A1(_1022_),
    .S(_1703_),
    .X(_1706_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(net668),
    .A1(_0982_),
    .S(_1702_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(net514),
    .A1(_1067_),
    .S(_1703_),
    .X(_1707_));
 sky130_fd_sc_hd__mux2_1 _5384_ (.A0(net515),
    .A1(_1030_),
    .S(_1702_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(net645),
    .A1(_1117_),
    .S(_1703_),
    .X(_1708_));
 sky130_fd_sc_hd__mux2_1 _5386_ (.A0(_1708_),
    .A1(_1075_),
    .S(_1702_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(net677),
    .A1(_1165_),
    .S(_1703_),
    .X(_1709_));
 sky130_fd_sc_hd__mux2_1 _5388_ (.A0(net678),
    .A1(_1125_),
    .S(_1702_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(net614),
    .A1(_1214_),
    .S(_1703_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(_1710_),
    .A1(_1172_),
    .S(_1702_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(net594),
    .A1(_1253_),
    .S(_1703_),
    .X(_1711_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(_1711_),
    .A1(_1219_),
    .S(_1702_),
    .X(_0249_));
 sky130_fd_sc_hd__or3b_4 _5393_ (.A(_0633_),
    .B(_0634_),
    .C_N(_1256_),
    .X(_1712_));
 sky130_fd_sc_hd__and3_4 _5394_ (.A(_0702_),
    .B(_0704_),
    .C(_1259_),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_1 _5395_ (.A0(net792),
    .A1(_0926_),
    .S(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(_0652_),
    .A1(net793),
    .S(_1712_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5397_ (.A0(net659),
    .A1(_0974_),
    .S(_1713_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(_0934_),
    .A1(_1715_),
    .S(_1712_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(net657),
    .A1(_1022_),
    .S(_1713_),
    .X(_1716_));
 sky130_fd_sc_hd__mux2_1 _5400_ (.A0(_0982_),
    .A1(net658),
    .S(_1712_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(net625),
    .A1(_1067_),
    .S(_1713_),
    .X(_1717_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(_1030_),
    .A1(net626),
    .S(_1712_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(net520),
    .A1(_1117_),
    .S(_1713_),
    .X(_1718_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(_1075_),
    .A1(_1718_),
    .S(_1712_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(net653),
    .A1(_1165_),
    .S(_1713_),
    .X(_1719_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(_1125_),
    .A1(net654),
    .S(_1712_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(net582),
    .A1(_1214_),
    .S(_1713_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(_1172_),
    .A1(_1720_),
    .S(_1712_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(net485),
    .A1(_1253_),
    .S(_1713_),
    .X(_1721_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(_1219_),
    .A1(_1721_),
    .S(_1712_),
    .X(_0257_));
 sky130_fd_sc_hd__or3_4 _5411_ (.A(net143),
    .B(net141),
    .C(net138),
    .X(_1722_));
 sky130_fd_sc_hd__or3_4 _5412_ (.A(net149),
    .B(net147),
    .C(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__a2111o_1 _5413_ (.A1(_3458_),
    .A2(net158),
    .B1(net156),
    .C1(net152),
    .D1(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__o41ai_2 _5414_ (.A1(net110),
    .A2(net155),
    .A3(net152),
    .A4(_1723_),
    .B1(\as1802.MHI[7] ),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2b_1 _5415_ (.A_N(\as1802.MHI[6] ),
    .B(net158),
    .Y(_1726_));
 sky130_fd_sc_hd__a21oi_1 _5416_ (.A1(\as1802.MHI[7] ),
    .A2(_1726_),
    .B1(net108),
    .Y(_1727_));
 sky130_fd_sc_hd__and2b_1 _5417_ (.A_N(_1726_),
    .B(_1725_),
    .X(_1728_));
 sky130_fd_sc_hd__nor2_1 _5418_ (.A(net152),
    .B(_1723_),
    .Y(_1729_));
 sky130_fd_sc_hd__or4_4 _5419_ (.A(net152),
    .B(net149),
    .C(net147),
    .D(_1722_),
    .X(_1730_));
 sky130_fd_sc_hd__o31a_1 _5420_ (.A1(net110),
    .A2(_1727_),
    .A3(_1730_),
    .B1(\as1802.MHI[6] ),
    .X(_1731_));
 sky130_fd_sc_hd__inv_2 _5421_ (.A(_1731_),
    .Y(_1732_));
 sky130_fd_sc_hd__a31oi_2 _5422_ (.A1(net156),
    .A2(_1726_),
    .A3(_1729_),
    .B1(_1725_),
    .Y(_1733_));
 sky130_fd_sc_hd__nor2_1 _5423_ (.A(net108),
    .B(_1731_),
    .Y(_1734_));
 sky130_fd_sc_hd__or2_4 _5424_ (.A(net108),
    .B(_1731_),
    .X(_1735_));
 sky130_fd_sc_hd__o311a_1 _5425_ (.A1(net110),
    .A2(net152),
    .A3(_1723_),
    .B1(net108),
    .C1(\as1802.MHI[6] ),
    .X(_1736_));
 sky130_fd_sc_hd__or2_1 _5426_ (.A(\as1802.MHI[5] ),
    .B(net110),
    .X(_1737_));
 sky130_fd_sc_hd__or2_4 _5427_ (.A(_1737_),
    .B(_1736_),
    .X(_1738_));
 sky130_fd_sc_hd__and3_1 _5428_ (.A(net107),
    .B(_1735_),
    .C(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__a31oi_4 _5429_ (.A1(net107),
    .A2(_1735_),
    .A3(_1738_),
    .B1(_1733_),
    .Y(_1740_));
 sky130_fd_sc_hd__a21oi_4 _5430_ (.A1(_1735_),
    .A2(_1738_),
    .B1(net107),
    .Y(_1741_));
 sky130_fd_sc_hd__or3_4 _5431_ (.A(_1723_),
    .B(_1740_),
    .C(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__nor2_1 _5432_ (.A(_1734_),
    .B(_1736_),
    .Y(_1743_));
 sky130_fd_sc_hd__xnor2_1 _5433_ (.A(_1737_),
    .B(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__mux2_4 _5434_ (.A0(_1744_),
    .A1(_1732_),
    .S(_1742_),
    .X(_1745_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(net152),
    .B(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(\as1802.MHI[5] ),
    .B(net110),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_1737_),
    .B(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__or4b_1 _5438_ (.A(_1723_),
    .B(_1740_),
    .C(_1741_),
    .D_N(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__o31ai_2 _5439_ (.A1(_1723_),
    .A2(_1740_),
    .A3(_1741_),
    .B1(\as1802.MHI[5] ),
    .Y(_1750_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_1749_),
    .B(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__and2_1 _5441_ (.A(net108),
    .B(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a21o_1 _5442_ (.A1(_1749_),
    .A2(_1750_),
    .B1(net156),
    .X(_1753_));
 sky130_fd_sc_hd__nor2_2 _5443_ (.A(\as1802.MHI[4] ),
    .B(net110),
    .Y(_1754_));
 sky130_fd_sc_hd__and3_1 _5444_ (.A(net156),
    .B(_1749_),
    .C(_1750_),
    .X(_1755_));
 sky130_fd_sc_hd__nor2_1 _5445_ (.A(_1752_),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__o21ai_1 _5446_ (.A1(_1754_),
    .A2(_1755_),
    .B1(_1753_),
    .Y(_1757_));
 sky130_fd_sc_hd__o221ai_4 _5447_ (.A1(net152),
    .A2(_1745_),
    .B1(_1754_),
    .B2(_1755_),
    .C1(_1753_),
    .Y(_1758_));
 sky130_fd_sc_hd__a21o_4 _5448_ (.A1(_1746_),
    .A2(_1758_),
    .B1(_3474_),
    .X(_1759_));
 sky130_fd_sc_hd__nor2_2 _5449_ (.A(net146),
    .B(_1722_),
    .Y(_1760_));
 sky130_fd_sc_hd__o21ai_2 _5450_ (.A1(_1739_),
    .A2(_1742_),
    .B1(_1733_),
    .Y(_1761_));
 sky130_fd_sc_hd__inv_2 _5451_ (.A(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__nand3_1 _5452_ (.A(_3474_),
    .B(_1746_),
    .C(_1758_),
    .Y(_1763_));
 sky130_fd_sc_hd__a31o_4 _5453_ (.A1(_3474_),
    .A2(_1746_),
    .A3(_1758_),
    .B1(_1762_),
    .X(_1764_));
 sky130_fd_sc_hd__nand3_4 _5454_ (.A(_1759_),
    .B(_1760_),
    .C(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__xnor2_1 _5455_ (.A(net107),
    .B(_1745_),
    .Y(_1766_));
 sky130_fd_sc_hd__xnor2_1 _5456_ (.A(_1757_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__mux2_2 _5457_ (.A0(_1767_),
    .A1(_1745_),
    .S(_1765_),
    .X(_1768_));
 sky130_fd_sc_hd__nor2_1 _5458_ (.A(net149),
    .B(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(net149),
    .B(_1768_),
    .Y(_1770_));
 sky130_fd_sc_hd__xnor2_1 _5460_ (.A(_1754_),
    .B(_1756_),
    .Y(_1771_));
 sky130_fd_sc_hd__a31o_1 _5461_ (.A1(_1759_),
    .A2(_1760_),
    .A3(_1764_),
    .B1(_1751_),
    .X(_1772_));
 sky130_fd_sc_hd__o21ai_1 _5462_ (.A1(_1765_),
    .A2(_1771_),
    .B1(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__o21a_1 _5463_ (.A1(_1765_),
    .A2(_1771_),
    .B1(_1772_),
    .X(_1774_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(net152),
    .B(_1773_),
    .Y(_1775_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_3473_),
    .B(_1774_),
    .Y(_1776_));
 sky130_fd_sc_hd__nor2_1 _5466_ (.A(_3459_),
    .B(net159),
    .Y(_1777_));
 sky130_fd_sc_hd__o2111ai_4 _5467_ (.A1(_1754_),
    .A2(_1777_),
    .B1(net255),
    .C1(_1760_),
    .D1(_1759_),
    .Y(_1778_));
 sky130_fd_sc_hd__a31o_4 _5468_ (.A1(_1759_),
    .A2(_1760_),
    .A3(_1764_),
    .B1(_3459_),
    .X(_1779_));
 sky130_fd_sc_hd__nand2_1 _5469_ (.A(_1778_),
    .B(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__a21oi_2 _5470_ (.A1(_1778_),
    .A2(_1779_),
    .B1(net155),
    .Y(_1781_));
 sky130_fd_sc_hd__nand3_2 _5471_ (.A(net155),
    .B(_1778_),
    .C(_1779_),
    .Y(_1782_));
 sky130_fd_sc_hd__and2b_1 _5472_ (.A_N(_1781_),
    .B(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__or2_2 _5473_ (.A(\as1802.MHI[3] ),
    .B(net110),
    .X(_1784_));
 sky130_fd_sc_hd__a21oi_1 _5474_ (.A1(_1782_),
    .A2(_1784_),
    .B1(_1781_),
    .Y(_1785_));
 sky130_fd_sc_hd__a221o_1 _5475_ (.A1(_3473_),
    .A2(_1774_),
    .B1(_1782_),
    .B2(_1784_),
    .C1(_1781_),
    .X(_1786_));
 sky130_fd_sc_hd__and2_1 _5476_ (.A(_1775_),
    .B(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__a31o_1 _5477_ (.A1(_1770_),
    .A2(_1775_),
    .A3(_1786_),
    .B1(_1769_),
    .X(_1788_));
 sky130_fd_sc_hd__a31o_1 _5478_ (.A1(_1759_),
    .A2(_1760_),
    .A3(_1763_),
    .B1(_1761_),
    .X(_1789_));
 sky130_fd_sc_hd__nand2_1 _5479_ (.A(net146),
    .B(_1761_),
    .Y(_1790_));
 sky130_fd_sc_hd__nor2_1 _5480_ (.A(net146),
    .B(_1789_),
    .Y(_1791_));
 sky130_fd_sc_hd__nand2_1 _5481_ (.A(\as1802.MHI[3] ),
    .B(net110),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_1775_),
    .B(_1776_),
    .Y(_1793_));
 sky130_fd_sc_hd__and2b_1 _5483_ (.A_N(_1769_),
    .B(_1770_),
    .X(_1794_));
 sky130_fd_sc_hd__a21oi_4 _5484_ (.A1(_1788_),
    .A2(_1790_),
    .B1(_1791_),
    .Y(_1795_));
 sky130_fd_sc_hd__nor2_4 _5485_ (.A(_1722_),
    .B(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__or4b_4 _5486_ (.A(net146),
    .B(net226),
    .C(_1789_),
    .D_N(_1788_),
    .X(_1797_));
 sky130_fd_sc_hd__o21a_1 _5487_ (.A1(_1789_),
    .A2(_1796_),
    .B1(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__or2_2 _5488_ (.A(net143),
    .B(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__xnor2_1 _5489_ (.A(_1787_),
    .B(_1794_),
    .Y(_1800_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(_1768_),
    .A1(_1800_),
    .S(_1796_),
    .X(_1801_));
 sky130_fd_sc_hd__or2_4 _5491_ (.A(net146),
    .B(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__nand2_1 _5492_ (.A(net146),
    .B(_1801_),
    .Y(_1803_));
 sky130_fd_sc_hd__nand2_1 _5493_ (.A(_1802_),
    .B(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__xnor2_1 _5494_ (.A(_1785_),
    .B(_1793_),
    .Y(_1805_));
 sky130_fd_sc_hd__mux2_4 _5495_ (.A0(_1773_),
    .A1(_1805_),
    .S(_1796_),
    .X(_1806_));
 sky130_fd_sc_hd__or2_4 _5496_ (.A(net149),
    .B(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__and2_4 _5497_ (.A(_1806_),
    .B(net149),
    .X(_1808_));
 sky130_fd_sc_hd__inv_2 _5498_ (.A(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__xor2_1 _5499_ (.A(_1783_),
    .B(_1784_),
    .X(_1810_));
 sky130_fd_sc_hd__or3_4 _5500_ (.A(_1722_),
    .B(_1795_),
    .C(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__o21ai_1 _5501_ (.A1(_1780_),
    .A2(_1796_),
    .B1(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__o21a_1 _5502_ (.A1(_1780_),
    .A2(_1796_),
    .B1(_1811_),
    .X(_1813_));
 sky130_fd_sc_hd__nor2_1 _5503_ (.A(net152),
    .B(_1812_),
    .Y(_1814_));
 sky130_fd_sc_hd__nor2_1 _5504_ (.A(_3473_),
    .B(_1813_),
    .Y(_1815_));
 sky130_fd_sc_hd__o21ai_2 _5505_ (.A1(net226),
    .A2(_1795_),
    .B1(\as1802.MHI[3] ),
    .Y(_1816_));
 sky130_fd_sc_hd__a211o_1 _5506_ (.A1(_1784_),
    .A2(_1792_),
    .B1(_1795_),
    .C1(net226),
    .X(_1817_));
 sky130_fd_sc_hd__and2_1 _5507_ (.A(_1816_),
    .B(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__a21o_1 _5508_ (.A1(_1816_),
    .A2(_1817_),
    .B1(net155),
    .X(_1819_));
 sky130_fd_sc_hd__nand2_1 _5509_ (.A(net155),
    .B(_1818_),
    .Y(_1820_));
 sky130_fd_sc_hd__nor2_1 _5510_ (.A(\as1802.MHI[2] ),
    .B(net111),
    .Y(_1821_));
 sky130_fd_sc_hd__a31o_1 _5511_ (.A1(net155),
    .A2(_1816_),
    .A3(_1817_),
    .B1(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__and2_1 _5512_ (.A(_1819_),
    .B(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__o2bb2a_2 _5513_ (.A1_N(_1819_),
    .A2_N(_1822_),
    .B1(_3473_),
    .B2(_1813_),
    .X(_1824_));
 sky130_fd_sc_hd__or2_1 _5514_ (.A(_1814_),
    .B(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__o21bai_4 _5515_ (.A1(_1814_),
    .A2(_1824_),
    .B1_N(_1808_),
    .Y(_1826_));
 sky130_fd_sc_hd__a21o_4 _5516_ (.A1(_1807_),
    .A2(_1826_),
    .B1(_1804_),
    .X(_1827_));
 sky130_fd_sc_hd__a211o_1 _5517_ (.A1(net143),
    .A2(_1798_),
    .B1(net138),
    .C1(net141),
    .X(_1828_));
 sky130_fd_sc_hd__a31oi_4 _5518_ (.A1(_1799_),
    .A2(_1802_),
    .A3(_1827_),
    .B1(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__a21oi_1 _5519_ (.A1(_1807_),
    .A2(_1809_),
    .B1(_1825_),
    .Y(_1830_));
 sky130_fd_sc_hd__and3_1 _5520_ (.A(_1807_),
    .B(_1809_),
    .C(_1825_),
    .X(_1831_));
 sky130_fd_sc_hd__or2_1 _5521_ (.A(_1830_),
    .B(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_4 _5522_ (.A0(_1806_),
    .A1(_1832_),
    .S(net248),
    .X(_1833_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(net146),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__or2_4 _5524_ (.A(net146),
    .B(_1833_),
    .X(_1835_));
 sky130_fd_sc_hd__inv_2 _5525_ (.A(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__or2_1 _5526_ (.A(_1814_),
    .B(_1815_),
    .X(_1837_));
 sky130_fd_sc_hd__xnor2_1 _5527_ (.A(_1823_),
    .B(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__mux2_2 _5528_ (.A0(_1812_),
    .A1(_1838_),
    .S(net248),
    .X(_1839_));
 sky130_fd_sc_hd__nor2_2 _5529_ (.A(net149),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__nand2_1 _5530_ (.A(_1819_),
    .B(_1820_),
    .Y(_1841_));
 sky130_fd_sc_hd__xnor2_1 _5531_ (.A(_1821_),
    .B(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__mux2_4 _5532_ (.A0(_1818_),
    .A1(_1842_),
    .S(net251),
    .X(_1843_));
 sky130_fd_sc_hd__nor2_4 _5533_ (.A(net152),
    .B(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__nand2_4 _5534_ (.A(_1843_),
    .B(net152),
    .Y(_1845_));
 sky130_fd_sc_hd__nor2_1 _5535_ (.A(_3460_),
    .B(net159),
    .Y(_1846_));
 sky130_fd_sc_hd__or2_1 _5536_ (.A(_1821_),
    .B(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__inv_2 _5537_ (.A(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__a311o_1 _5538_ (.A1(_1799_),
    .A2(_1802_),
    .A3(_1827_),
    .B1(_1828_),
    .C1(_1847_),
    .X(_1849_));
 sky130_fd_sc_hd__a311o_1 _5539_ (.A1(_1799_),
    .A2(_1802_),
    .A3(_1827_),
    .B1(_1828_),
    .C1(_1848_),
    .X(_1850_));
 sky130_fd_sc_hd__o21a_1 _5540_ (.A1(\as1802.MHI[2] ),
    .A2(net219),
    .B1(_1849_),
    .X(_1851_));
 sky130_fd_sc_hd__o211ai_1 _5541_ (.A1(\as1802.MHI[2] ),
    .A2(net237),
    .B1(_1849_),
    .C1(net108),
    .Y(_1852_));
 sky130_fd_sc_hd__nor2_1 _5542_ (.A(\as1802.MHI[1] ),
    .B(net111),
    .Y(_1853_));
 sky130_fd_sc_hd__o211a_1 _5543_ (.A1(_3460_),
    .A2(net219),
    .B1(_1850_),
    .C1(net155),
    .X(_1854_));
 sky130_fd_sc_hd__o21ai_2 _5544_ (.A1(_1853_),
    .A2(_1854_),
    .B1(_1852_),
    .Y(_1855_));
 sky130_fd_sc_hd__a21o_1 _5545_ (.A1(_1845_),
    .A2(_1855_),
    .B1(_1844_),
    .X(_1856_));
 sky130_fd_sc_hd__nand2_1 _5546_ (.A(net149),
    .B(_1839_),
    .Y(_1857_));
 sky130_fd_sc_hd__a21oi_1 _5547_ (.A1(net223),
    .A2(_1857_),
    .B1(_1840_),
    .Y(_1858_));
 sky130_fd_sc_hd__a211o_4 _5548_ (.A1(_1856_),
    .A2(_1857_),
    .B1(_1836_),
    .C1(_1840_),
    .X(_1859_));
 sky130_fd_sc_hd__nand2_1 _5549_ (.A(_1834_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__a21o_1 _5550_ (.A1(_1802_),
    .A2(_1827_),
    .B1(net226),
    .X(_1861_));
 sky130_fd_sc_hd__a21o_1 _5551_ (.A1(net219),
    .A2(_1861_),
    .B1(_1798_),
    .X(_1862_));
 sky130_fd_sc_hd__xnor2_1 _5552_ (.A(net141),
    .B(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand3_1 _5553_ (.A(_1804_),
    .B(_1807_),
    .C(_1826_),
    .Y(_1864_));
 sky130_fd_sc_hd__nand2_1 _5554_ (.A(_1827_),
    .B(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__mux2_4 _5555_ (.A0(_1801_),
    .A1(_1865_),
    .S(net247),
    .X(_1866_));
 sky130_fd_sc_hd__xnor2_2 _5556_ (.A(net143),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__nor2_2 _5557_ (.A(_1863_),
    .B(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__a211o_1 _5558_ (.A1(net141),
    .A2(_1862_),
    .B1(_1866_),
    .C1(net143),
    .X(_1869_));
 sky130_fd_sc_hd__o21ai_2 _5559_ (.A1(net141),
    .A2(_1862_),
    .B1(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__a31oi_4 _5560_ (.A1(_1834_),
    .A2(_1859_),
    .A3(_1868_),
    .B1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__a31o_1 _5561_ (.A1(_1834_),
    .A2(net246),
    .A3(net253),
    .B1(_1870_),
    .X(_1872_));
 sky130_fd_sc_hd__nor2_4 _5562_ (.A(net138),
    .B(_1871_),
    .Y(_1873_));
 sky130_fd_sc_hd__xnor2_1 _5563_ (.A(_1860_),
    .B(_1867_),
    .Y(_1874_));
 sky130_fd_sc_hd__mux2_2 _5564_ (.A0(_1866_),
    .A1(_1874_),
    .S(_1873_),
    .X(_1875_));
 sky130_fd_sc_hd__xnor2_2 _5565_ (.A(net141),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__and2_1 _5566_ (.A(net138),
    .B(_1862_),
    .X(_1877_));
 sky130_fd_sc_hd__o21a_1 _5567_ (.A1(_1862_),
    .A2(_1873_),
    .B1(_1797_),
    .X(_1878_));
 sky130_fd_sc_hd__nor2_1 _5568_ (.A(net138),
    .B(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__or2_1 _5569_ (.A(_1876_),
    .B(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__nor3_1 _5570_ (.A(_1876_),
    .B(_1877_),
    .C(_1879_),
    .Y(_1881_));
 sky130_fd_sc_hd__or2_2 _5571_ (.A(_1877_),
    .B(_1880_),
    .X(_1882_));
 sky130_fd_sc_hd__and2b_1 _5572_ (.A_N(_1840_),
    .B(_1857_),
    .X(_1883_));
 sky130_fd_sc_hd__xnor2_1 _5573_ (.A(net224),
    .B(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__mux2_2 _5574_ (.A0(_1839_),
    .A1(_1884_),
    .S(_1873_),
    .X(_1885_));
 sky130_fd_sc_hd__or2_1 _5575_ (.A(net146),
    .B(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__xnor2_2 _5576_ (.A(net148),
    .B(_1885_),
    .Y(_1887_));
 sky130_fd_sc_hd__nand2_1 _5577_ (.A(_1834_),
    .B(net254),
    .Y(_1888_));
 sky130_fd_sc_hd__xnor2_1 _5578_ (.A(_1858_),
    .B(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(_1833_),
    .A1(_1889_),
    .S(_1873_),
    .X(_1890_));
 sky130_fd_sc_hd__xnor2_1 _5580_ (.A(net250),
    .B(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__nor2_1 _5581_ (.A(_1887_),
    .B(_1891_),
    .Y(_1892_));
 sky130_fd_sc_hd__or2_1 _5582_ (.A(_1887_),
    .B(_1891_),
    .X(_1893_));
 sky130_fd_sc_hd__and2b_1 _5583_ (.A_N(_1844_),
    .B(_1845_),
    .X(_1894_));
 sky130_fd_sc_hd__nor2_1 _5584_ (.A(net249),
    .B(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__and2_1 _5585_ (.A(_1855_),
    .B(_1894_),
    .X(_1896_));
 sky130_fd_sc_hd__a21o_1 _5586_ (.A1(_3478_),
    .A2(net240),
    .B1(_1843_),
    .X(_1897_));
 sky130_fd_sc_hd__or4_4 _5587_ (.A(net138),
    .B(_1871_),
    .C(_1895_),
    .D(_1896_),
    .X(_1898_));
 sky130_fd_sc_hd__and2_1 _5588_ (.A(_1897_),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__and3_1 _5589_ (.A(net149),
    .B(_1897_),
    .C(_1898_),
    .X(_1900_));
 sky130_fd_sc_hd__xnor2_1 _5590_ (.A(net108),
    .B(_1851_),
    .Y(_1901_));
 sky130_fd_sc_hd__or3b_4 _5591_ (.A(net138),
    .B(_1871_),
    .C_N(_1853_),
    .X(_1902_));
 sky130_fd_sc_hd__a21o_1 _5592_ (.A1(_3478_),
    .A2(_1872_),
    .B1(net108),
    .X(_1903_));
 sky130_fd_sc_hd__a21o_1 _5593_ (.A1(_1902_),
    .A2(_1903_),
    .B1(_1901_),
    .X(_1904_));
 sky130_fd_sc_hd__nand3_2 _5594_ (.A(_1901_),
    .B(_1902_),
    .C(_1903_),
    .Y(_1905_));
 sky130_fd_sc_hd__and2_1 _5595_ (.A(_1904_),
    .B(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__a21oi_1 _5596_ (.A1(_1904_),
    .A2(_1905_),
    .B1(net152),
    .Y(_1907_));
 sky130_fd_sc_hd__a21o_1 _5597_ (.A1(_1904_),
    .A2(_1905_),
    .B1(net152),
    .X(_1908_));
 sky130_fd_sc_hd__and3_1 _5598_ (.A(net154),
    .B(_1904_),
    .C(_1905_),
    .X(_1909_));
 sky130_fd_sc_hd__or2_1 _5599_ (.A(_1907_),
    .B(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__a31o_1 _5600_ (.A1(net159),
    .A2(_3478_),
    .A3(_1872_),
    .B1(_3461_),
    .X(_1911_));
 sky130_fd_sc_hd__and2_1 _5601_ (.A(_1902_),
    .B(net239),
    .X(_1912_));
 sky130_fd_sc_hd__a21oi_1 _5602_ (.A1(_1902_),
    .A2(net239),
    .B1(net155),
    .Y(_1913_));
 sky130_fd_sc_hd__a21o_1 _5603_ (.A1(_1902_),
    .A2(_1911_),
    .B1(net155),
    .X(_1914_));
 sky130_fd_sc_hd__nand2_1 _5604_ (.A(_3462_),
    .B(net159),
    .Y(_1915_));
 sky130_fd_sc_hd__and3_1 _5605_ (.A(net155),
    .B(_1902_),
    .C(_1911_),
    .X(_1916_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(\as1802.MHI[0] ),
    .B(net111),
    .Y(_1917_));
 sky130_fd_sc_hd__nand2_1 _5607_ (.A(_1915_),
    .B(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__inv_2 _5608_ (.A(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__or2_1 _5609_ (.A(_1913_),
    .B(net889),
    .X(_1920_));
 sky130_fd_sc_hd__a31o_1 _5610_ (.A1(_3462_),
    .A2(net159),
    .A3(_1914_),
    .B1(net889),
    .X(_1921_));
 sky130_fd_sc_hd__a21oi_1 _5611_ (.A1(_1897_),
    .A2(net241),
    .B1(net149),
    .Y(_1922_));
 sky130_fd_sc_hd__or2_1 _5612_ (.A(net150),
    .B(_1899_),
    .X(_1923_));
 sky130_fd_sc_hd__o211a_1 _5613_ (.A1(_1909_),
    .A2(_1921_),
    .B1(_1923_),
    .C1(_1908_),
    .X(_1924_));
 sky130_fd_sc_hd__nor2_1 _5614_ (.A(net221),
    .B(_1922_),
    .Y(_1925_));
 sky130_fd_sc_hd__nor4b_1 _5615_ (.A(_1907_),
    .B(_1909_),
    .C(_1920_),
    .D_N(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__a211o_1 _5616_ (.A1(_1904_),
    .A2(_1905_),
    .B1(net154),
    .C1(net220),
    .X(_1927_));
 sky130_fd_sc_hd__a2111o_1 _5617_ (.A1(_1914_),
    .A2(_1917_),
    .B1(_1922_),
    .C1(_1916_),
    .D1(_1900_),
    .X(_1928_));
 sky130_fd_sc_hd__o311a_1 _5618_ (.A1(_1907_),
    .A2(_1909_),
    .A3(_1928_),
    .B1(_1927_),
    .C1(_1923_),
    .X(_1929_));
 sky130_fd_sc_hd__or2_1 _5619_ (.A(net221),
    .B(_1924_),
    .X(_1930_));
 sky130_fd_sc_hd__or3_4 _5620_ (.A(_1893_),
    .B(net221),
    .C(_1924_),
    .X(_1931_));
 sky130_fd_sc_hd__nand4_1 _5621_ (.A(_1881_),
    .B(_1892_),
    .C(_1919_),
    .D(_1926_),
    .Y(_1932_));
 sky130_fd_sc_hd__or3b_4 _5622_ (.A(_1929_),
    .B(_1893_),
    .C_N(_1881_),
    .X(_1933_));
 sky130_fd_sc_hd__a211o_1 _5623_ (.A1(net250),
    .A2(_1890_),
    .B1(_1885_),
    .C1(net148),
    .X(_1934_));
 sky130_fd_sc_hd__o21a_1 _5624_ (.A1(net144),
    .A2(_1890_),
    .B1(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__o32a_1 _5625_ (.A1(net141),
    .A2(_1875_),
    .A3(_1877_),
    .B1(_1878_),
    .B2(net138),
    .X(_1936_));
 sky130_fd_sc_hd__o31a_2 _5626_ (.A1(_1877_),
    .A2(_1880_),
    .A3(_1935_),
    .B1(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__o21ai_4 _5627_ (.A1(_1882_),
    .A2(_1931_),
    .B1(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__a22o_1 _5628_ (.A1(net131),
    .A2(net150),
    .B1(net147),
    .B2(net134),
    .X(_1939_));
 sky130_fd_sc_hd__inv_2 _5629_ (.A(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__and4_1 _5630_ (.A(net131),
    .B(net134),
    .C(net150),
    .D(net147),
    .X(_1941_));
 sky130_fd_sc_hd__and4b_1 _5631_ (.A_N(_1941_),
    .B(net153),
    .C(net129),
    .D(_1939_),
    .X(_1942_));
 sky130_fd_sc_hd__o22a_1 _5632_ (.A1(_3435_),
    .A2(net107),
    .B1(_1940_),
    .B2(_1941_),
    .X(_1943_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(net135),
    .B(net245),
    .Y(_1944_));
 sky130_fd_sc_hd__or3_1 _5634_ (.A(_1942_),
    .B(_1943_),
    .C(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(net128),
    .B(net153),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_2 _5636_ (.A(net129),
    .B(net150),
    .Y(_1947_));
 sky130_fd_sc_hd__o21a_1 _5637_ (.A1(_3436_),
    .A2(_3475_),
    .B1(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__and4_1 _5638_ (.A(net129),
    .B(net131),
    .C(net150),
    .D(net147),
    .X(_1949_));
 sky130_fd_sc_hd__nor2_1 _5639_ (.A(_1948_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__xnor2_1 _5640_ (.A(_1946_),
    .B(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__a22o_1 _5641_ (.A1(net134),
    .A2(net244),
    .B1(net141),
    .B2(net135),
    .X(_1952_));
 sky130_fd_sc_hd__inv_2 _5642_ (.A(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__and4_1 _5643_ (.A(net134),
    .B(net135),
    .C(net244),
    .D(net140),
    .X(_1954_));
 sky130_fd_sc_hd__or3b_1 _5644_ (.A(_1953_),
    .B(_1954_),
    .C_N(_1951_),
    .X(_1955_));
 sky130_fd_sc_hd__o21bai_1 _5645_ (.A1(_1953_),
    .A2(_1954_),
    .B1_N(_1951_),
    .Y(_1956_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_1955_),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__or2_1 _5647_ (.A(_1945_),
    .B(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__nand2_1 _5648_ (.A(net122),
    .B(net158),
    .Y(_1959_));
 sky130_fd_sc_hd__o211a_1 _5649_ (.A1(_1941_),
    .A2(_1942_),
    .B1(net124),
    .C1(net156),
    .X(_1960_));
 sky130_fd_sc_hd__a211oi_1 _5650_ (.A1(net124),
    .A2(net156),
    .B1(_1941_),
    .C1(_1942_),
    .Y(_1961_));
 sky130_fd_sc_hd__nor2_1 _5651_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__xnor2_1 _5652_ (.A(_1959_),
    .B(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(_1945_),
    .B(_1957_),
    .Y(_1964_));
 sky130_fd_sc_hd__and2_1 _5654_ (.A(_1958_),
    .B(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__nand2_1 _5655_ (.A(_1963_),
    .B(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__nand2_1 _5656_ (.A(net122),
    .B(net155),
    .Y(_1967_));
 sky130_fd_sc_hd__a31o_1 _5657_ (.A1(net128),
    .A2(net153),
    .A3(_1950_),
    .B1(_1949_),
    .X(_1968_));
 sky130_fd_sc_hd__and3_1 _5658_ (.A(net122),
    .B(net155),
    .C(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__xnor2_1 _5659_ (.A(_1967_),
    .B(_1968_),
    .Y(_1970_));
 sky130_fd_sc_hd__and3_1 _5660_ (.A(net120),
    .B(net159),
    .C(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__a21oi_1 _5661_ (.A1(net120),
    .A2(net159),
    .B1(_1970_),
    .Y(_1972_));
 sky130_fd_sc_hd__nor2_1 _5662_ (.A(_1971_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__a22o_1 _5663_ (.A1(net128),
    .A2(net150),
    .B1(net148),
    .B2(net129),
    .X(_1974_));
 sky130_fd_sc_hd__inv_2 _5664_ (.A(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__and4_1 _5665_ (.A(net128),
    .B(net130),
    .C(net149),
    .D(net148),
    .X(_1976_));
 sky130_fd_sc_hd__and4b_1 _5666_ (.A_N(_1976_),
    .B(net152),
    .C(net125),
    .D(_1974_),
    .X(_1977_));
 sky130_fd_sc_hd__o2bb2a_1 _5667_ (.A1_N(net124),
    .A2_N(net152),
    .B1(_1975_),
    .B2(_1976_),
    .X(_1978_));
 sky130_fd_sc_hd__a22o_1 _5668_ (.A1(net134),
    .A2(net140),
    .B1(net137),
    .B2(net136),
    .X(_1979_));
 sky130_fd_sc_hd__inv_2 _5669_ (.A(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__and4_1 _5670_ (.A(net134),
    .B(net136),
    .C(net140),
    .D(net137),
    .X(_1981_));
 sky130_fd_sc_hd__and4b_1 _5671_ (.A_N(_1981_),
    .B(net144),
    .C(net131),
    .D(_1979_),
    .X(_1982_));
 sky130_fd_sc_hd__o22a_1 _5672_ (.A1(_3436_),
    .A2(_3476_),
    .B1(_1980_),
    .B2(_1981_),
    .X(_1983_));
 sky130_fd_sc_hd__nor2_1 _5673_ (.A(_1982_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__nand2_1 _5674_ (.A(_1954_),
    .B(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__or2_1 _5675_ (.A(_1954_),
    .B(_1984_),
    .X(_1986_));
 sky130_fd_sc_hd__nand2_1 _5676_ (.A(_1985_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__or3_1 _5677_ (.A(_1977_),
    .B(_1978_),
    .C(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__o21ai_1 _5678_ (.A1(_1977_),
    .A2(_1978_),
    .B1(_1987_),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _5679_ (.A(_1988_),
    .B(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__nor2_2 _5680_ (.A(_1955_),
    .B(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__and2_1 _5681_ (.A(_1955_),
    .B(_1990_),
    .X(_1992_));
 sky130_fd_sc_hd__nor2_1 _5682_ (.A(_1991_),
    .B(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__and2_2 _5683_ (.A(_1973_),
    .B(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__nor2_1 _5684_ (.A(_1973_),
    .B(_1993_),
    .Y(_1995_));
 sky130_fd_sc_hd__a211oi_2 _5685_ (.A1(_1958_),
    .A2(_1966_),
    .B1(_1994_),
    .C1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__a31o_1 _5686_ (.A1(net122),
    .A2(net158),
    .A3(_1962_),
    .B1(_1960_),
    .X(_1997_));
 sky130_fd_sc_hd__o211a_1 _5687_ (.A1(_1994_),
    .A2(_1995_),
    .B1(_1958_),
    .C1(_1966_),
    .X(_1998_));
 sky130_fd_sc_hd__nor2_1 _5688_ (.A(_1996_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__and2_1 _5689_ (.A(_1997_),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__o211a_1 _5690_ (.A1(_1976_),
    .A2(_1977_),
    .B1(net121),
    .C1(net156),
    .X(_2001_));
 sky130_fd_sc_hd__inv_2 _5691_ (.A(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__a211o_1 _5692_ (.A1(net121),
    .A2(net156),
    .B1(_1976_),
    .C1(_1977_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _5693_ (.A(_2002_),
    .B(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__nor2_2 _5694_ (.A(_3434_),
    .B(_3475_),
    .Y(_2005_));
 sky130_fd_sc_hd__a21oi_1 _5695_ (.A1(net124),
    .A2(net150),
    .B1(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__and3_1 _5696_ (.A(net125),
    .B(net150),
    .C(_2005_),
    .X(_2007_));
 sky130_fd_sc_hd__nor2_1 _5697_ (.A(_2006_),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__and3_1 _5698_ (.A(net122),
    .B(net153),
    .C(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__a21oi_1 _5699_ (.A1(net122),
    .A2(net153),
    .B1(_2008_),
    .Y(_2010_));
 sky130_fd_sc_hd__nor2_1 _5700_ (.A(_2009_),
    .B(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__or2_1 _5701_ (.A(_1981_),
    .B(_1982_),
    .X(_2012_));
 sky130_fd_sc_hd__a22o_1 _5702_ (.A1(net131),
    .A2(net140),
    .B1(net137),
    .B2(net134),
    .X(_2013_));
 sky130_fd_sc_hd__inv_2 _5703_ (.A(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__and4_1 _5704_ (.A(net131),
    .B(net134),
    .C(net140),
    .D(net137),
    .X(_2015_));
 sky130_fd_sc_hd__and4b_1 _5705_ (.A_N(_2015_),
    .B(net245),
    .C(net129),
    .D(_2013_),
    .X(_2016_));
 sky130_fd_sc_hd__o22a_1 _5706_ (.A1(_3435_),
    .A2(_3476_),
    .B1(_2014_),
    .B2(_2015_),
    .X(_2017_));
 sky130_fd_sc_hd__nor2_1 _5707_ (.A(_2016_),
    .B(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(_2012_),
    .B(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__xor2_1 _5709_ (.A(_2012_),
    .B(_2018_),
    .X(_2020_));
 sky130_fd_sc_hd__nand2_1 _5710_ (.A(_2011_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__or2_1 _5711_ (.A(_2011_),
    .B(_2020_),
    .X(_2022_));
 sky130_fd_sc_hd__nand2_1 _5712_ (.A(_2021_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__a21oi_1 _5713_ (.A1(_1985_),
    .A2(_1988_),
    .B1(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__and3_1 _5714_ (.A(_1985_),
    .B(_1988_),
    .C(_2023_),
    .X(_2025_));
 sky130_fd_sc_hd__or3_2 _5715_ (.A(_2004_),
    .B(_2024_),
    .C(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__o21ai_2 _5716_ (.A1(_2024_),
    .A2(_2025_),
    .B1(_2004_),
    .Y(_2027_));
 sky130_fd_sc_hd__o211ai_4 _5717_ (.A1(_1991_),
    .A2(_1994_),
    .B1(_2026_),
    .C1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__a211o_1 _5718_ (.A1(_2026_),
    .A2(_2027_),
    .B1(_1991_),
    .C1(_1994_),
    .X(_2029_));
 sky130_fd_sc_hd__o211ai_4 _5719_ (.A1(_1969_),
    .A2(_1971_),
    .B1(_2028_),
    .C1(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__a211o_1 _5720_ (.A1(_2028_),
    .A2(_2029_),
    .B1(_1969_),
    .C1(_1971_),
    .X(_2031_));
 sky130_fd_sc_hd__o211ai_2 _5721_ (.A1(_1996_),
    .A2(_2000_),
    .B1(_2030_),
    .C1(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__a211o_1 _5722_ (.A1(_2030_),
    .A2(_2031_),
    .B1(_1996_),
    .C1(_2000_),
    .X(_2033_));
 sky130_fd_sc_hd__and2_1 _5723_ (.A(_2032_),
    .B(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__and4_1 _5724_ (.A(net134),
    .B(net136),
    .C(net151),
    .D(net148),
    .X(_2035_));
 sky130_fd_sc_hd__nand2_2 _5725_ (.A(net131),
    .B(net154),
    .Y(_2036_));
 sky130_fd_sc_hd__o22a_1 _5726_ (.A1(_3437_),
    .A2(net106),
    .B1(_3475_),
    .B2(_3438_),
    .X(_2037_));
 sky130_fd_sc_hd__or2_1 _5727_ (.A(_2035_),
    .B(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nor2_1 _5728_ (.A(_2036_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__o211a_1 _5729_ (.A1(_2035_),
    .A2(_2039_),
    .B1(net127),
    .C1(net157),
    .X(_2040_));
 sky130_fd_sc_hd__a211oi_1 _5730_ (.A1(net127),
    .A2(net157),
    .B1(_2035_),
    .C1(_2039_),
    .Y(_2041_));
 sky130_fd_sc_hd__nor2_1 _5731_ (.A(_2040_),
    .B(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__and3_1 _5732_ (.A(net124),
    .B(net158),
    .C(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__a21oi_1 _5733_ (.A1(net124),
    .A2(net158),
    .B1(_2042_),
    .Y(_2044_));
 sky130_fd_sc_hd__nor2_1 _5734_ (.A(_2043_),
    .B(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__o21ai_1 _5735_ (.A1(_1942_),
    .A2(_1943_),
    .B1(_1944_),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _5736_ (.A(_1945_),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__inv_2 _5737_ (.A(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_2045_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__or2_1 _5739_ (.A(_1963_),
    .B(_1965_),
    .X(_2050_));
 sky130_fd_sc_hd__nand2_1 _5740_ (.A(_1966_),
    .B(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__or2_1 _5741_ (.A(_2049_),
    .B(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__nand2_1 _5742_ (.A(_2049_),
    .B(_2051_),
    .Y(_2053_));
 sky130_fd_sc_hd__and2_1 _5743_ (.A(_2052_),
    .B(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__o21ai_2 _5744_ (.A1(_2040_),
    .A2(_2043_),
    .B1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__xnor2_2 _5745_ (.A(_1997_),
    .B(_1999_),
    .Y(_2056_));
 sky130_fd_sc_hd__a21oi_2 _5746_ (.A1(_2052_),
    .A2(_2055_),
    .B1(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__and3_1 _5747_ (.A(_2052_),
    .B(_2055_),
    .C(_2056_),
    .X(_2058_));
 sky130_fd_sc_hd__and2_1 _5748_ (.A(_2036_),
    .B(_2038_),
    .X(_2059_));
 sky130_fd_sc_hd__nor2_1 _5749_ (.A(_2039_),
    .B(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__and4_1 _5750_ (.A(net134),
    .B(net136),
    .C(net154),
    .D(net151),
    .X(_2061_));
 sky130_fd_sc_hd__a21oi_1 _5751_ (.A1(net129),
    .A2(net157),
    .B1(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__and3_1 _5752_ (.A(net129),
    .B(net157),
    .C(_2061_),
    .X(_2063_));
 sky130_fd_sc_hd__and4bb_1 _5753_ (.A_N(_2062_),
    .B_N(_2063_),
    .C(net128),
    .D(net158),
    .X(_2064_));
 sky130_fd_sc_hd__o22a_1 _5754_ (.A1(_3434_),
    .A2(net111),
    .B1(_2062_),
    .B2(_2063_),
    .X(_2065_));
 sky130_fd_sc_hd__nor2_1 _5755_ (.A(_2064_),
    .B(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(_2060_),
    .B(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__or2_1 _5757_ (.A(_2045_),
    .B(_2048_),
    .X(_2068_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_2049_),
    .B(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__or2_1 _5759_ (.A(_2067_),
    .B(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(_2067_),
    .B(_2069_),
    .Y(_2071_));
 sky130_fd_sc_hd__and2_1 _5761_ (.A(_2070_),
    .B(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__o21ai_1 _5762_ (.A1(_2063_),
    .A2(_2064_),
    .B1(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__or3_1 _5763_ (.A(_2040_),
    .B(_2043_),
    .C(_2054_),
    .X(_2074_));
 sky130_fd_sc_hd__nand2_1 _5764_ (.A(_2055_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__a21o_1 _5765_ (.A1(_2070_),
    .A2(_2073_),
    .B1(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__or3_1 _5766_ (.A(_2063_),
    .B(_2064_),
    .C(_2072_),
    .X(_2077_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_2073_),
    .B(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__or2_1 _5768_ (.A(_2060_),
    .B(_2066_),
    .X(_2079_));
 sky130_fd_sc_hd__and2_1 _5769_ (.A(_2067_),
    .B(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__and4_1 _5770_ (.A(net129),
    .B(net131),
    .C(net158),
    .D(net156),
    .X(_2081_));
 sky130_fd_sc_hd__or4_1 _5771_ (.A(_3435_),
    .B(_3436_),
    .C(net110),
    .D(net109),
    .X(_2082_));
 sky130_fd_sc_hd__a22o_1 _5772_ (.A1(net129),
    .A2(net158),
    .B1(net156),
    .B2(net131),
    .X(_2083_));
 sky130_fd_sc_hd__o22a_1 _5773_ (.A1(_3437_),
    .A2(net107),
    .B1(net106),
    .B2(_3438_),
    .X(_2084_));
 sky130_fd_sc_hd__nor2_1 _5774_ (.A(_2061_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__and3_1 _5775_ (.A(_2082_),
    .B(_2083_),
    .C(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__o21ai_1 _5776_ (.A1(_2081_),
    .A2(_2086_),
    .B1(_2080_),
    .Y(_2087_));
 sky130_fd_sc_hd__or3_1 _5777_ (.A(_2080_),
    .B(_2081_),
    .C(_2086_),
    .X(_2088_));
 sky130_fd_sc_hd__and2_1 _5778_ (.A(_2087_),
    .B(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__a21o_1 _5779_ (.A1(_2082_),
    .A2(_2083_),
    .B1(_2085_),
    .X(_2090_));
 sky130_fd_sc_hd__and2b_1 _5780_ (.A_N(_2086_),
    .B(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__nand2_2 _5781_ (.A(net133),
    .B(net157),
    .Y(_2092_));
 sky130_fd_sc_hd__and4_1 _5782_ (.A(net131),
    .B(net134),
    .C(net160),
    .D(net157),
    .X(_2093_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(net136),
    .B(net154),
    .Y(_2094_));
 sky130_fd_sc_hd__o21ai_2 _5784_ (.A1(_3436_),
    .A2(net111),
    .B1(_2092_),
    .Y(_2095_));
 sky130_fd_sc_hd__and2b_1 _5785_ (.A_N(_2093_),
    .B(_2095_),
    .X(_2096_));
 sky130_fd_sc_hd__a31o_1 _5786_ (.A1(net136),
    .A2(net154),
    .A3(_2095_),
    .B1(_2093_),
    .X(_2097_));
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(net134),
    .B(net160),
    .Y(_2098_));
 sky130_fd_sc_hd__and4_1 _5788_ (.A(net134),
    .B(net136),
    .C(net158),
    .D(net156),
    .X(_2099_));
 sky130_fd_sc_hd__inv_2 _5789_ (.A(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__xnor2_1 _5790_ (.A(_2094_),
    .B(_2096_),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(_2099_),
    .B(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__xnor2_1 _5792_ (.A(_2091_),
    .B(_2097_),
    .Y(_2103_));
 sky130_fd_sc_hd__or2_1 _5793_ (.A(_2102_),
    .B(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__a21boi_1 _5794_ (.A1(_2091_),
    .A2(_2097_),
    .B1_N(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__nand2b_1 _5795_ (.A_N(_2105_),
    .B(_2089_),
    .Y(_2106_));
 sky130_fd_sc_hd__a21oi_2 _5796_ (.A1(_2087_),
    .A2(_2106_),
    .B1(_2078_),
    .Y(_2107_));
 sky130_fd_sc_hd__nand3_1 _5797_ (.A(_2070_),
    .B(_2073_),
    .C(_2075_),
    .Y(_2108_));
 sky130_fd_sc_hd__nand3_2 _5798_ (.A(_2076_),
    .B(_2107_),
    .C(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__a211oi_2 _5799_ (.A1(_2076_),
    .A2(_2109_),
    .B1(_2057_),
    .C1(_2058_),
    .Y(_2110_));
 sky130_fd_sc_hd__or3_1 _5800_ (.A(_2034_),
    .B(_2057_),
    .C(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__o21ai_1 _5801_ (.A1(_2057_),
    .A2(_2110_),
    .B1(_2034_),
    .Y(_2112_));
 sky130_fd_sc_hd__and3_1 _5802_ (.A(_3510_),
    .B(_2111_),
    .C(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__a21o_1 _5803_ (.A1(net97),
    .A2(net229),
    .B1(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__or4_1 _5804_ (.A(_3553_),
    .B(_0542_),
    .C(_0574_),
    .D(_0592_),
    .X(_2115_));
 sky130_fd_sc_hd__or3b_1 _5805_ (.A(net170),
    .B(net171),
    .C_N(net168),
    .X(_2116_));
 sky130_fd_sc_hd__o22a_1 _5806_ (.A1(_0510_),
    .A2(_0528_),
    .B1(_2116_),
    .B2(net119),
    .X(_2117_));
 sky130_fd_sc_hd__a21o_1 _5807_ (.A1(net162),
    .A2(_3498_),
    .B1(_3494_),
    .X(_2118_));
 sky130_fd_sc_hd__nor2_1 _5808_ (.A(_3486_),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__nor4_1 _5809_ (.A(_3501_),
    .B(_2115_),
    .C(_2117_),
    .D(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__or4_4 _5810_ (.A(_3501_),
    .B(_2115_),
    .C(_2117_),
    .D(_2119_),
    .X(_2121_));
 sky130_fd_sc_hd__nor2_2 _5811_ (.A(_3489_),
    .B(_3576_),
    .Y(_2122_));
 sky130_fd_sc_hd__a221o_1 _5812_ (.A1(_3489_),
    .A2(_2114_),
    .B1(_2122_),
    .B2(net135),
    .C1(_2121_),
    .X(_2123_));
 sky130_fd_sc_hd__o211a_1 _5813_ (.A1(net294),
    .A2(net79),
    .B1(_2123_),
    .C1(net212),
    .X(_0258_));
 sky130_fd_sc_hd__and2b_1 _5814_ (.A_N(_2024_),
    .B(_2026_),
    .X(_2124_));
 sky130_fd_sc_hd__a22o_1 _5815_ (.A1(net122),
    .A2(net149),
    .B1(net147),
    .B2(net124),
    .X(_2125_));
 sky130_fd_sc_hd__and4_1 _5816_ (.A(net122),
    .B(net124),
    .C(net149),
    .D(net147),
    .X(_2126_));
 sky130_fd_sc_hd__nand4_1 _5817_ (.A(net122),
    .B(net125),
    .C(net149),
    .D(net147),
    .Y(_2127_));
 sky130_fd_sc_hd__and4_1 _5818_ (.A(net121),
    .B(net152),
    .C(_2125_),
    .D(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__o2bb2a_1 _5819_ (.A1_N(_2125_),
    .A2_N(_2127_),
    .B1(_3433_),
    .B2(_3473_),
    .X(_2129_));
 sky130_fd_sc_hd__nor2_1 _5820_ (.A(_2128_),
    .B(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__or2_1 _5821_ (.A(_2015_),
    .B(_2016_),
    .X(_2131_));
 sky130_fd_sc_hd__a22o_1 _5822_ (.A1(net129),
    .A2(net140),
    .B1(net137),
    .B2(net131),
    .X(_2132_));
 sky130_fd_sc_hd__inv_2 _5823_ (.A(_2132_),
    .Y(_2133_));
 sky130_fd_sc_hd__and4_1 _5824_ (.A(net129),
    .B(net131),
    .C(net140),
    .D(net137),
    .X(_2134_));
 sky130_fd_sc_hd__and4b_1 _5825_ (.A_N(_2134_),
    .B(net242),
    .C(net128),
    .D(_2132_),
    .X(_2135_));
 sky130_fd_sc_hd__o22a_1 _5826_ (.A1(_3434_),
    .A2(_3476_),
    .B1(_2133_),
    .B2(_2134_),
    .X(_2136_));
 sky130_fd_sc_hd__nor2_1 _5827_ (.A(_2135_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_2131_),
    .B(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__xor2_1 _5829_ (.A(_2131_),
    .B(_2137_),
    .X(_2139_));
 sky130_fd_sc_hd__nand2_1 _5830_ (.A(_2130_),
    .B(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__or2_1 _5831_ (.A(_2130_),
    .B(_2139_),
    .X(_2141_));
 sky130_fd_sc_hd__nand2_1 _5832_ (.A(_2140_),
    .B(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__a21o_1 _5833_ (.A1(_2019_),
    .A2(_2021_),
    .B1(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__nand3_1 _5834_ (.A(_2019_),
    .B(_2021_),
    .C(_2142_),
    .Y(_2144_));
 sky130_fd_sc_hd__o211ai_1 _5835_ (.A1(_2007_),
    .A2(_2009_),
    .B1(_2143_),
    .C1(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__a211o_1 _5836_ (.A1(_2143_),
    .A2(_2144_),
    .B1(_2007_),
    .C1(_2009_),
    .X(_2146_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_2145_),
    .B(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__xnor2_1 _5838_ (.A(_2124_),
    .B(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__or2_1 _5839_ (.A(_2002_),
    .B(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__nand2_1 _5840_ (.A(_2002_),
    .B(_2148_),
    .Y(_2150_));
 sky130_fd_sc_hd__nand2_1 _5841_ (.A(_2149_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__a21o_1 _5842_ (.A1(_2028_),
    .A2(_2030_),
    .B1(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__and3_1 _5843_ (.A(_2028_),
    .B(_2030_),
    .C(_2151_),
    .X(_2153_));
 sky130_fd_sc_hd__inv_2 _5844_ (.A(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__nand2_1 _5845_ (.A(_2152_),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__a21o_1 _5846_ (.A1(_2032_),
    .A2(_2112_),
    .B1(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__a31oi_1 _5847_ (.A1(_2032_),
    .A2(_2112_),
    .A3(_2155_),
    .B1(net97),
    .Y(_2157_));
 sky130_fd_sc_hd__a22o_1 _5848_ (.A1(net97),
    .A2(_1873_),
    .B1(_2156_),
    .B2(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__a221o_1 _5849_ (.A1(net134),
    .A2(_2122_),
    .B1(_2158_),
    .B2(_3489_),
    .C1(_2121_),
    .X(_2159_));
 sky130_fd_sc_hd__o211a_1 _5850_ (.A1(net300),
    .A2(net79),
    .B1(_2159_),
    .C1(net212),
    .X(_0259_));
 sky130_fd_sc_hd__o21ai_1 _5851_ (.A1(_2124_),
    .A2(_2147_),
    .B1(_2149_),
    .Y(_2160_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_2143_),
    .B(_2145_),
    .Y(_2161_));
 sky130_fd_sc_hd__a22oi_1 _5853_ (.A1(net121),
    .A2(net149),
    .B1(net147),
    .B2(net123),
    .Y(_2162_));
 sky130_fd_sc_hd__and4_1 _5854_ (.A(net121),
    .B(net123),
    .C(net149),
    .D(net147),
    .X(_2163_));
 sky130_fd_sc_hd__nor2_1 _5855_ (.A(_2162_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__or2_1 _5856_ (.A(_2134_),
    .B(_2135_),
    .X(_2165_));
 sky130_fd_sc_hd__nand2_4 _5857_ (.A(net124),
    .B(net145),
    .Y(_2166_));
 sky130_fd_sc_hd__a22o_1 _5858_ (.A1(net127),
    .A2(net140),
    .B1(net137),
    .B2(net129),
    .X(_2167_));
 sky130_fd_sc_hd__inv_2 _5859_ (.A(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__and4_1 _5860_ (.A(net127),
    .B(net129),
    .C(net140),
    .D(net137),
    .X(_2169_));
 sky130_fd_sc_hd__nor2_1 _5861_ (.A(_2168_),
    .B(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__xnor2_1 _5862_ (.A(_2166_),
    .B(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__and2_1 _5863_ (.A(_2165_),
    .B(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__xor2_1 _5864_ (.A(_2165_),
    .B(_2171_),
    .X(_2173_));
 sky130_fd_sc_hd__and2_1 _5865_ (.A(_2164_),
    .B(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__nor2_1 _5866_ (.A(_2164_),
    .B(_2173_),
    .Y(_2175_));
 sky130_fd_sc_hd__or2_1 _5867_ (.A(_2174_),
    .B(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__a21o_1 _5868_ (.A1(_2138_),
    .A2(_2140_),
    .B1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nand3_1 _5869_ (.A(_2138_),
    .B(_2140_),
    .C(_2176_),
    .Y(_2178_));
 sky130_fd_sc_hd__o211ai_2 _5870_ (.A1(_2126_),
    .A2(_2128_),
    .B1(_2177_),
    .C1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__a211o_1 _5871_ (.A1(_2177_),
    .A2(_2178_),
    .B1(_2126_),
    .C1(_2128_),
    .X(_2180_));
 sky130_fd_sc_hd__and3_1 _5872_ (.A(_2161_),
    .B(_2179_),
    .C(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__a21oi_1 _5873_ (.A1(_2179_),
    .A2(_2180_),
    .B1(_2161_),
    .Y(_2182_));
 sky130_fd_sc_hd__nor2_1 _5874_ (.A(_2181_),
    .B(_2182_),
    .Y(_2183_));
 sky130_fd_sc_hd__and2_1 _5875_ (.A(_2160_),
    .B(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__xnor2_1 _5876_ (.A(_2160_),
    .B(_2183_),
    .Y(_2185_));
 sky130_fd_sc_hd__and3_1 _5877_ (.A(_2152_),
    .B(_2156_),
    .C(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__a21oi_1 _5878_ (.A1(_2152_),
    .A2(_2156_),
    .B1(_2185_),
    .Y(_2187_));
 sky130_fd_sc_hd__or2_1 _5879_ (.A(net97),
    .B(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__o2bb2a_1 _5880_ (.A1_N(net97),
    .A2_N(net219),
    .B1(_2186_),
    .B2(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__nor2_1 _5881_ (.A(_3488_),
    .B(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__a21o_1 _5882_ (.A1(net131),
    .A2(_2122_),
    .B1(_2121_),
    .X(_2191_));
 sky130_fd_sc_hd__o221a_1 _5883_ (.A1(net726),
    .A2(net79),
    .B1(_2190_),
    .B2(_2191_),
    .C1(net212),
    .X(_0260_));
 sky130_fd_sc_hd__a31o_1 _5884_ (.A1(net124),
    .A2(net242),
    .A3(_2167_),
    .B1(_2169_),
    .X(_2192_));
 sky130_fd_sc_hd__o2bb2a_1 _5885_ (.A1_N(net124),
    .A2_N(net140),
    .B1(_3478_),
    .B2(_3434_),
    .X(_2193_));
 sky130_fd_sc_hd__and4_1 _5886_ (.A(net124),
    .B(net128),
    .C(net140),
    .D(net137),
    .X(_2194_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(_2193_),
    .B(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__and3_1 _5888_ (.A(net122),
    .B(net242),
    .C(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__a21oi_1 _5889_ (.A1(net122),
    .A2(net242),
    .B1(_2195_),
    .Y(_2197_));
 sky130_fd_sc_hd__nor2_1 _5890_ (.A(_2196_),
    .B(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__and2_1 _5891_ (.A(_2192_),
    .B(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__nor2_1 _5892_ (.A(_2192_),
    .B(_2198_),
    .Y(_2200_));
 sky130_fd_sc_hd__nor2_1 _5893_ (.A(_2199_),
    .B(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__and3_1 _5894_ (.A(net121),
    .B(net147),
    .C(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__a21oi_1 _5895_ (.A1(net121),
    .A2(net147),
    .B1(_2201_),
    .Y(_2203_));
 sky130_fd_sc_hd__nor2_1 _5896_ (.A(_2202_),
    .B(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__o21a_1 _5897_ (.A1(_2172_),
    .A2(_2174_),
    .B1(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__nor3_1 _5898_ (.A(_2172_),
    .B(_2174_),
    .C(_2204_),
    .Y(_2206_));
 sky130_fd_sc_hd__nor2_1 _5899_ (.A(_2205_),
    .B(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__and2_1 _5900_ (.A(_2163_),
    .B(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__nor2_1 _5901_ (.A(_2163_),
    .B(_2207_),
    .Y(_2209_));
 sky130_fd_sc_hd__or2_1 _5902_ (.A(_2208_),
    .B(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__a21o_1 _5903_ (.A1(_2177_),
    .A2(_2179_),
    .B1(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__nand3_1 _5904_ (.A(_2177_),
    .B(_2179_),
    .C(_2210_),
    .Y(_2212_));
 sky130_fd_sc_hd__and3_1 _5905_ (.A(_2181_),
    .B(_2211_),
    .C(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__a21oi_1 _5906_ (.A1(_2211_),
    .A2(_2212_),
    .B1(_2181_),
    .Y(_2214_));
 sky130_fd_sc_hd__nor2_1 _5907_ (.A(_2213_),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__o21a_1 _5908_ (.A1(_2184_),
    .A2(_2187_),
    .B1(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__o31ai_1 _5909_ (.A1(_2184_),
    .A2(_2187_),
    .A3(_2215_),
    .B1(_3510_),
    .Y(_2217_));
 sky130_fd_sc_hd__a2bb2o_1 _5910_ (.A1_N(_2216_),
    .A2_N(_2217_),
    .B1(net98),
    .B2(_1796_),
    .X(_2218_));
 sky130_fd_sc_hd__a221o_1 _5911_ (.A1(net130),
    .A2(_2122_),
    .B1(_2218_),
    .B2(_3489_),
    .C1(_2121_),
    .X(_2219_));
 sky130_fd_sc_hd__o211a_1 _5912_ (.A1(net304),
    .A2(net79),
    .B1(_2219_),
    .C1(net213),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_1 _5913_ (.A(_2194_),
    .B(_2196_),
    .Y(_2220_));
 sky130_fd_sc_hd__and2_1 _5914_ (.A(net123),
    .B(net142),
    .X(_2221_));
 sky130_fd_sc_hd__nand2_1 _5915_ (.A(net123),
    .B(net142),
    .Y(_2222_));
 sky130_fd_sc_hd__a21oi_1 _5916_ (.A1(net124),
    .A2(net139),
    .B1(_2221_),
    .Y(_2223_));
 sky130_fd_sc_hd__and3_1 _5917_ (.A(net124),
    .B(net139),
    .C(_2221_),
    .X(_2224_));
 sky130_fd_sc_hd__and4bb_1 _5918_ (.A_N(_2223_),
    .B_N(_2224_),
    .C(net121),
    .D(net242),
    .X(_2225_));
 sky130_fd_sc_hd__o22a_1 _5919_ (.A1(_3433_),
    .A2(_3476_),
    .B1(_2223_),
    .B2(_2224_),
    .X(_2226_));
 sky130_fd_sc_hd__nor2_1 _5920_ (.A(_2225_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__o21a_1 _5921_ (.A1(_2194_),
    .A2(_2196_),
    .B1(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__xnor2_1 _5922_ (.A(_2220_),
    .B(_2227_),
    .Y(_2229_));
 sky130_fd_sc_hd__nor3_1 _5923_ (.A(_2199_),
    .B(_2202_),
    .C(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__o21a_1 _5924_ (.A1(_2199_),
    .A2(_2202_),
    .B1(_2229_),
    .X(_2231_));
 sky130_fd_sc_hd__nor2_1 _5925_ (.A(_2230_),
    .B(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__o21ai_1 _5926_ (.A1(_2205_),
    .A2(_2208_),
    .B1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__or3_1 _5927_ (.A(_2205_),
    .B(_2208_),
    .C(_2232_),
    .X(_2234_));
 sky130_fd_sc_hd__nand2_1 _5928_ (.A(_2233_),
    .B(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__nor2_1 _5929_ (.A(_2211_),
    .B(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__and2_1 _5930_ (.A(_2211_),
    .B(_2235_),
    .X(_2237_));
 sky130_fd_sc_hd__nor2_1 _5931_ (.A(_2236_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__o21a_1 _5932_ (.A1(_2213_),
    .A2(_2216_),
    .B1(_2238_),
    .X(_2239_));
 sky130_fd_sc_hd__nor3_1 _5933_ (.A(_2213_),
    .B(_2216_),
    .C(_2238_),
    .Y(_2240_));
 sky130_fd_sc_hd__o21ai_1 _5934_ (.A1(_2239_),
    .A2(_2240_),
    .B1(_3510_),
    .Y(_2241_));
 sky130_fd_sc_hd__a21oi_1 _5935_ (.A1(net98),
    .A2(_1765_),
    .B1(_3488_),
    .Y(_2242_));
 sky130_fd_sc_hd__a221o_1 _5936_ (.A1(net127),
    .A2(_2122_),
    .B1(_2241_),
    .B2(_2242_),
    .C1(_2121_),
    .X(_2243_));
 sky130_fd_sc_hd__o211a_1 _5937_ (.A1(net308),
    .A2(net79),
    .B1(_2243_),
    .C1(net213),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(net120),
    .B(net142),
    .Y(_2244_));
 sky130_fd_sc_hd__nand2_1 _5939_ (.A(net123),
    .B(net139),
    .Y(_2245_));
 sky130_fd_sc_hd__xor2_1 _5940_ (.A(_2244_),
    .B(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__or3_1 _5941_ (.A(_2224_),
    .B(_2225_),
    .C(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__o21ai_1 _5942_ (.A1(_2224_),
    .A2(_2225_),
    .B1(_2246_),
    .Y(_2248_));
 sky130_fd_sc_hd__and2_1 _5943_ (.A(_2247_),
    .B(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__or2_1 _5944_ (.A(_2228_),
    .B(_2231_),
    .X(_2250_));
 sky130_fd_sc_hd__xnor2_1 _5945_ (.A(_2249_),
    .B(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__nor2_1 _5946_ (.A(_2233_),
    .B(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__and2_1 _5947_ (.A(_2233_),
    .B(_2251_),
    .X(_2253_));
 sky130_fd_sc_hd__nor2_1 _5948_ (.A(_2252_),
    .B(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__o21a_1 _5949_ (.A1(_2236_),
    .A2(_2239_),
    .B1(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__o31ai_1 _5950_ (.A1(_2236_),
    .A2(_2239_),
    .A3(_2254_),
    .B1(_3510_),
    .Y(_2256_));
 sky130_fd_sc_hd__o22a_1 _5951_ (.A1(_3510_),
    .A2(_1742_),
    .B1(_2255_),
    .B2(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__nor2_1 _5952_ (.A(_3488_),
    .B(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__a21o_1 _5953_ (.A1(net125),
    .A2(_2122_),
    .B1(_2121_),
    .X(_2259_));
 sky130_fd_sc_hd__o221a_1 _5954_ (.A1(net319),
    .A2(net79),
    .B1(_2258_),
    .B2(_2259_),
    .C1(net213),
    .X(_0263_));
 sky130_fd_sc_hd__or4_1 _5955_ (.A(_3510_),
    .B(_1727_),
    .C(_1728_),
    .D(_1730_),
    .X(_2260_));
 sky130_fd_sc_hd__and2_1 _5956_ (.A(_2228_),
    .B(_2249_),
    .X(_2261_));
 sky130_fd_sc_hd__nand2_2 _5957_ (.A(net120),
    .B(net139),
    .Y(_2262_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_2222_),
    .B(_2248_),
    .Y(_2263_));
 sky130_fd_sc_hd__mux2_1 _5959_ (.A0(_2263_),
    .A1(_2248_),
    .S(_2262_),
    .X(_2264_));
 sky130_fd_sc_hd__xnor2_1 _5960_ (.A(_2261_),
    .B(_2264_),
    .Y(_2265_));
 sky130_fd_sc_hd__and3_1 _5961_ (.A(_2231_),
    .B(_2249_),
    .C(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__a21oi_1 _5962_ (.A1(_2231_),
    .A2(_2249_),
    .B1(_2265_),
    .Y(_2267_));
 sky130_fd_sc_hd__nor2_1 _5963_ (.A(_2266_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__nor3_1 _5964_ (.A(_2252_),
    .B(_2255_),
    .C(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__o21a_1 _5965_ (.A1(_2252_),
    .A2(_2255_),
    .B1(_2268_),
    .X(_2270_));
 sky130_fd_sc_hd__o31ai_1 _5966_ (.A1(net98),
    .A2(_2269_),
    .A3(_2270_),
    .B1(_2260_),
    .Y(_2271_));
 sky130_fd_sc_hd__a221o_1 _5967_ (.A1(net122),
    .A2(_2122_),
    .B1(_2271_),
    .B2(_3489_),
    .C1(_2121_),
    .X(_2272_));
 sky130_fd_sc_hd__o211a_1 _5968_ (.A1(net296),
    .A2(net79),
    .B1(_2272_),
    .C1(net213),
    .X(_0264_));
 sky130_fd_sc_hd__o21ba_1 _5969_ (.A1(_2261_),
    .A2(_2263_),
    .B1_N(_2262_),
    .X(_2273_));
 sky130_fd_sc_hd__or4_1 _5970_ (.A(net98),
    .B(_2266_),
    .C(_2270_),
    .D(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__a21oi_1 _5971_ (.A1(net98),
    .A2(_1724_),
    .B1(_3488_),
    .Y(_2275_));
 sky130_fd_sc_hd__a221o_1 _5972_ (.A1(net121),
    .A2(_2122_),
    .B1(_2274_),
    .B2(_2275_),
    .C1(_2121_),
    .X(_2276_));
 sky130_fd_sc_hd__o211a_1 _5973_ (.A1(net375),
    .A2(net79),
    .B1(_2276_),
    .C1(net213),
    .X(_0265_));
 sky130_fd_sc_hd__or4_1 _5974_ (.A(net173),
    .B(_3440_),
    .C(_0498_),
    .D(_0521_),
    .X(_2277_));
 sky130_fd_sc_hd__a211o_1 _5975_ (.A1(net171),
    .A2(_0508_),
    .B1(_3528_),
    .C1(net173),
    .X(_2278_));
 sky130_fd_sc_hd__inv_2 _5976_ (.A(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__or4_1 _5977_ (.A(net172),
    .B(_3440_),
    .C(net171),
    .D(_3522_),
    .X(_2280_));
 sky130_fd_sc_hd__nor2_1 _5978_ (.A(net824),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__nor2_1 _5979_ (.A(_0534_),
    .B(_0581_),
    .Y(_2282_));
 sky130_fd_sc_hd__nand2_1 _5980_ (.A(_3432_),
    .B(_0526_),
    .Y(_2283_));
 sky130_fd_sc_hd__o2111a_1 _5981_ (.A1(net164),
    .A2(_0514_),
    .B1(_0526_),
    .C1(_3578_),
    .D1(_3432_),
    .X(_2284_));
 sky130_fd_sc_hd__a2111oi_1 _5982_ (.A1(_3432_),
    .A2(_3498_),
    .B1(_2281_),
    .C1(_2282_),
    .D1(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__a31o_1 _5983_ (.A1(_2277_),
    .A2(_2278_),
    .A3(_2285_),
    .B1(net102),
    .X(_2286_));
 sky130_fd_sc_hd__o32a_1 _5984_ (.A1(_3440_),
    .A2(_3553_),
    .A3(_0543_),
    .B1(_0544_),
    .B2(_0560_),
    .X(_2287_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_3496_),
    .B(_3506_),
    .Y(_2288_));
 sky130_fd_sc_hd__a31o_1 _5986_ (.A1(_0524_),
    .A2(_0666_),
    .A3(_2288_),
    .B1(_0560_),
    .X(_2289_));
 sky130_fd_sc_hd__o21a_1 _5987_ (.A1(net172),
    .A2(_0533_),
    .B1(_0679_),
    .X(_2290_));
 sky130_fd_sc_hd__or3b_1 _5988_ (.A(net163),
    .B(_3531_),
    .C_N(_3576_),
    .X(_2291_));
 sky130_fd_sc_hd__a2111o_1 _5989_ (.A1(_3432_),
    .A2(_2291_),
    .B1(_3541_),
    .C1(_3537_),
    .D1(net102),
    .X(_2292_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(net104),
    .B(_0678_),
    .Y(_2293_));
 sky130_fd_sc_hd__a32o_1 _5991_ (.A1(net104),
    .A2(_3579_),
    .A3(_0678_),
    .B1(_0578_),
    .B2(_3552_),
    .X(_2294_));
 sky130_fd_sc_hd__a31o_1 _5992_ (.A1(_3539_),
    .A2(_3540_),
    .A3(_0576_),
    .B1(net102),
    .X(_2295_));
 sky130_fd_sc_hd__o211a_1 _5993_ (.A1(_0539_),
    .A2(_2290_),
    .B1(_2295_),
    .C1(_0562_),
    .X(_2296_));
 sky130_fd_sc_hd__and4b_1 _5994_ (.A_N(_2294_),
    .B(_2296_),
    .C(_2289_),
    .D(_2292_),
    .X(_2297_));
 sky130_fd_sc_hd__nand4_2 _5995_ (.A(net209),
    .B(_2286_),
    .C(_2287_),
    .D(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__xor2_1 _5996_ (.A(net331),
    .B(net280),
    .X(_2299_));
 sky130_fd_sc_hd__a221o_1 _5997_ (.A1(net377),
    .A2(_3447_),
    .B1(net369),
    .B2(_3449_),
    .C1(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__xor2_1 _5998_ (.A(net333),
    .B(net292),
    .X(_2301_));
 sky130_fd_sc_hd__xor2_1 _5999_ (.A(net340),
    .B(net286),
    .X(_2302_));
 sky130_fd_sc_hd__a22o_1 _6000_ (.A1(_3446_),
    .A2(net306),
    .B1(net373),
    .B2(_3451_),
    .X(_2303_));
 sky130_fd_sc_hd__a221o_1 _6001_ (.A1(_3448_),
    .A2(net298),
    .B1(_3450_),
    .B2(net282),
    .C1(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__a221o_1 _6002_ (.A1(net461),
    .A2(_3453_),
    .B1(net371),
    .B2(_3455_),
    .C1(_2301_),
    .X(_2305_));
 sky130_fd_sc_hd__a221o_1 _6003_ (.A1(_3452_),
    .A2(net302),
    .B1(_3454_),
    .B2(net290),
    .C1(_2302_),
    .X(_2306_));
 sky130_fd_sc_hd__or4_4 _6004_ (.A(_2300_),
    .B(_2304_),
    .C(_2305_),
    .D(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__o21ba_1 _6005_ (.A1(_3551_),
    .A2(_2307_),
    .B1_N(_3546_),
    .X(_2308_));
 sky130_fd_sc_hd__o21a_1 _6006_ (.A1(net366),
    .A2(_2308_),
    .B1(net352),
    .X(_2309_));
 sky130_fd_sc_hd__nor2_1 _6007_ (.A(_2298_),
    .B(net367),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_4 _6008_ (.A(_3457_),
    .B(_2307_),
    .Y(_2310_));
 sky130_fd_sc_hd__a221oi_1 _6009_ (.A1(_3457_),
    .A2(_3548_),
    .B1(_2310_),
    .B2(net352),
    .C1(_2298_),
    .Y(_0267_));
 sky130_fd_sc_hd__a21oi_1 _6010_ (.A1(_3547_),
    .A2(_2310_),
    .B1(_3555_),
    .Y(_2311_));
 sky130_fd_sc_hd__nor2_1 _6011_ (.A(_3464_),
    .B(_2311_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_1 _6012_ (.A1(_0557_),
    .A2(_0666_),
    .B1(_2277_),
    .Y(_2312_));
 sky130_fd_sc_hd__or3b_1 _6013_ (.A(_2312_),
    .B(_2281_),
    .C_N(_0582_),
    .X(_2313_));
 sky130_fd_sc_hd__o21a_1 _6014_ (.A1(_0524_),
    .A2(_0557_),
    .B1(net104),
    .X(_2314_));
 sky130_fd_sc_hd__and4_1 _6015_ (.A(net209),
    .B(_3539_),
    .C(_3540_),
    .D(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__a21oi_1 _6016_ (.A1(_0533_),
    .A2(_2291_),
    .B1(net172),
    .Y(_2316_));
 sky130_fd_sc_hd__o32a_1 _6017_ (.A1(net172),
    .A2(_3485_),
    .A3(_3492_),
    .B1(_0557_),
    .B2(_2288_),
    .X(_2317_));
 sky130_fd_sc_hd__a21oi_1 _6018_ (.A1(_3499_),
    .A2(_3525_),
    .B1(net172),
    .Y(_2318_));
 sky130_fd_sc_hd__or4b_1 _6019_ (.A(_0575_),
    .B(_2318_),
    .C(_2316_),
    .D_N(_2317_),
    .X(_2319_));
 sky130_fd_sc_hd__or4b_1 _6020_ (.A(_2282_),
    .B(_2319_),
    .C(_2284_),
    .D_N(_2315_),
    .X(_2320_));
 sky130_fd_sc_hd__or3_2 _6021_ (.A(_2279_),
    .B(_2313_),
    .C(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__nor2_2 _6022_ (.A(net174),
    .B(_3527_),
    .Y(_2322_));
 sky130_fd_sc_hd__mux2_1 _6023_ (.A0(_3465_),
    .A1(_0889_),
    .S(_0584_),
    .X(_2323_));
 sky130_fd_sc_hd__o21a_1 _6024_ (.A1(net166),
    .A2(_0889_),
    .B1(_1335_),
    .X(_2324_));
 sky130_fd_sc_hd__a21oi_4 _6025_ (.A1(net95),
    .A2(_0513_),
    .B1(_0516_),
    .Y(_2325_));
 sky130_fd_sc_hd__o21a_1 _6026_ (.A1(\as1802.instr_latch[7] ),
    .A2(_3493_),
    .B1(_3524_),
    .X(_2326_));
 sky130_fd_sc_hd__inv_2 _6027_ (.A(net87),
    .Y(_2327_));
 sky130_fd_sc_hd__o211a_1 _6028_ (.A1(net95),
    .A2(_0799_),
    .B1(net87),
    .C1(_3528_),
    .X(_2328_));
 sky130_fd_sc_hd__o221a_1 _6029_ (.A1(net94),
    .A2(_2323_),
    .B1(_2324_),
    .B2(_2325_),
    .C1(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__a21oi_1 _6030_ (.A1(_0420_),
    .A2(_2327_),
    .B1(_2329_),
    .Y(_2330_));
 sky130_fd_sc_hd__o22a_1 _6031_ (.A1(_0800_),
    .A2(_2322_),
    .B1(_2330_),
    .B2(\as1802.instr_cycle[0] ),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _6032_ (.A0(_2331_),
    .A1(net272),
    .S(net77),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _6033_ (.A0(_0729_),
    .A1(_0880_),
    .S(net118),
    .X(_2332_));
 sky130_fd_sc_hd__inv_2 _6034_ (.A(_2332_),
    .Y(_2333_));
 sky130_fd_sc_hd__nor2_1 _6035_ (.A(net93),
    .B(_0880_),
    .Y(_2334_));
 sky130_fd_sc_hd__a211o_1 _6036_ (.A1(\as1802.regs[2][1] ),
    .A2(net93),
    .B1(_2334_),
    .C1(net94),
    .X(_2335_));
 sky130_fd_sc_hd__o21a_1 _6037_ (.A1(_2325_),
    .A2(_2333_),
    .B1(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__o221a_1 _6038_ (.A1(net95),
    .A2(_0730_),
    .B1(_2336_),
    .B2(net96),
    .C1(net87),
    .X(_2337_));
 sky130_fd_sc_hd__nor2_1 _6039_ (.A(_0428_),
    .B(net87),
    .Y(_2338_));
 sky130_fd_sc_hd__o32a_1 _6040_ (.A1(net173),
    .A2(_2337_),
    .A3(_2338_),
    .B1(_0730_),
    .B2(net88),
    .X(_2339_));
 sky130_fd_sc_hd__mux2_1 _6041_ (.A0(_2339_),
    .A1(net268),
    .S(net77),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _6042_ (.A0(_0738_),
    .A1(_0871_),
    .S(net118),
    .X(_2340_));
 sky130_fd_sc_hd__inv_2 _6043_ (.A(_2340_),
    .Y(_2341_));
 sky130_fd_sc_hd__nor2_1 _6044_ (.A(net91),
    .B(_0871_),
    .Y(_2342_));
 sky130_fd_sc_hd__a211o_1 _6045_ (.A1(\as1802.regs[2][2] ),
    .A2(net91),
    .B1(_2342_),
    .C1(net94),
    .X(_2343_));
 sky130_fd_sc_hd__o21a_1 _6046_ (.A1(_2325_),
    .A2(_2341_),
    .B1(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__o221a_1 _6047_ (.A1(net95),
    .A2(_0739_),
    .B1(_2344_),
    .B2(net96),
    .C1(net87),
    .X(_2345_));
 sky130_fd_sc_hd__nor2_1 _6048_ (.A(_0412_),
    .B(net87),
    .Y(_2346_));
 sky130_fd_sc_hd__o32a_1 _6049_ (.A1(net172),
    .A2(_2345_),
    .A3(_2346_),
    .B1(_0739_),
    .B2(net88),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _6050_ (.A0(_2347_),
    .A1(net266),
    .S(net77),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _6051_ (.A0(_0748_),
    .A1(_0860_),
    .S(net118),
    .X(_2348_));
 sky130_fd_sc_hd__inv_2 _6052_ (.A(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__nor2_1 _6053_ (.A(net91),
    .B(_0860_),
    .Y(_2350_));
 sky130_fd_sc_hd__a211o_1 _6054_ (.A1(\as1802.regs[2][3] ),
    .A2(net91),
    .B1(_2350_),
    .C1(net94),
    .X(_2351_));
 sky130_fd_sc_hd__o21a_1 _6055_ (.A1(_2325_),
    .A2(_2349_),
    .B1(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__o221a_1 _6056_ (.A1(net95),
    .A2(_0749_),
    .B1(_2352_),
    .B2(net96),
    .C1(net87),
    .X(_2353_));
 sky130_fd_sc_hd__nor2_1 _6057_ (.A(_0404_),
    .B(net87),
    .Y(_2354_));
 sky130_fd_sc_hd__o32a_1 _6058_ (.A1(net173),
    .A2(_2353_),
    .A3(_2354_),
    .B1(_0749_),
    .B2(net88),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _6059_ (.A0(_2355_),
    .A1(net264),
    .S(net77),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _6060_ (.A0(_0758_),
    .A1(_0849_),
    .S(net118),
    .X(_2356_));
 sky130_fd_sc_hd__inv_2 _6061_ (.A(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(net91),
    .B(_0849_),
    .Y(_2358_));
 sky130_fd_sc_hd__a211o_1 _6063_ (.A1(\as1802.regs[2][4] ),
    .A2(net91),
    .B1(_2358_),
    .C1(net94),
    .X(_2359_));
 sky130_fd_sc_hd__o21a_1 _6064_ (.A1(_2325_),
    .A2(_2357_),
    .B1(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__o221a_1 _6065_ (.A1(net95),
    .A2(_0759_),
    .B1(_2360_),
    .B2(net96),
    .C1(net87),
    .X(_2361_));
 sky130_fd_sc_hd__nor2_1 _6066_ (.A(_0396_),
    .B(net87),
    .Y(_2362_));
 sky130_fd_sc_hd__o32a_1 _6067_ (.A1(net173),
    .A2(_2361_),
    .A3(_2362_),
    .B1(_0759_),
    .B2(net88),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _6068_ (.A0(_2363_),
    .A1(net262),
    .S(net77),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _6069_ (.A0(_0768_),
    .A1(_0840_),
    .S(net117),
    .X(_2364_));
 sky130_fd_sc_hd__inv_2 _6070_ (.A(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__nor2_1 _6071_ (.A(net91),
    .B(_0840_),
    .Y(_2366_));
 sky130_fd_sc_hd__a211o_1 _6072_ (.A1(\as1802.regs[2][5] ),
    .A2(net93),
    .B1(_2366_),
    .C1(net94),
    .X(_2367_));
 sky130_fd_sc_hd__o21a_1 _6073_ (.A1(_2325_),
    .A2(_2365_),
    .B1(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__o221a_1 _6074_ (.A1(net95),
    .A2(_0769_),
    .B1(_2368_),
    .B2(net96),
    .C1(net87),
    .X(_2369_));
 sky130_fd_sc_hd__nor2_1 _6075_ (.A(_0388_),
    .B(net87),
    .Y(_2370_));
 sky130_fd_sc_hd__o32a_1 _6076_ (.A1(net174),
    .A2(_2369_),
    .A3(_2370_),
    .B1(_0769_),
    .B2(net88),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _6077_ (.A0(_2371_),
    .A1(net256),
    .S(net77),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _6078_ (.A0(_0778_),
    .A1(_0905_),
    .S(net118),
    .X(_2372_));
 sky130_fd_sc_hd__inv_2 _6079_ (.A(_2372_),
    .Y(_2373_));
 sky130_fd_sc_hd__nor2_1 _6080_ (.A(net92),
    .B(_0905_),
    .Y(_2374_));
 sky130_fd_sc_hd__a211o_1 _6081_ (.A1(\as1802.regs[2][6] ),
    .A2(net92),
    .B1(_2374_),
    .C1(net94),
    .X(_2375_));
 sky130_fd_sc_hd__o21a_1 _6082_ (.A1(_2325_),
    .A2(_2373_),
    .B1(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__o221a_1 _6083_ (.A1(net95),
    .A2(_0779_),
    .B1(_2376_),
    .B2(net96),
    .C1(net86),
    .X(_2377_));
 sky130_fd_sc_hd__nor2_1 _6084_ (.A(_0441_),
    .B(net86),
    .Y(_2378_));
 sky130_fd_sc_hd__o32a_1 _6085_ (.A1(net174),
    .A2(_2377_),
    .A3(_2378_),
    .B1(_0779_),
    .B2(net88),
    .X(_2379_));
 sky130_fd_sc_hd__mux2_1 _6086_ (.A0(_2379_),
    .A1(net258),
    .S(_2321_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _6087_ (.A0(_0788_),
    .A1(_0916_),
    .S(net118),
    .X(_2380_));
 sky130_fd_sc_hd__inv_2 _6088_ (.A(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__nor2_1 _6089_ (.A(net92),
    .B(_0916_),
    .Y(_2382_));
 sky130_fd_sc_hd__a211o_1 _6090_ (.A1(\as1802.regs[2][7] ),
    .A2(net92),
    .B1(_2382_),
    .C1(net94),
    .X(_2383_));
 sky130_fd_sc_hd__o21a_1 _6091_ (.A1(_2325_),
    .A2(_2381_),
    .B1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__o221a_1 _6092_ (.A1(net95),
    .A2(_0789_),
    .B1(_2384_),
    .B2(net96),
    .C1(net86),
    .X(_2385_));
 sky130_fd_sc_hd__nor2_1 _6093_ (.A(_0451_),
    .B(net86),
    .Y(_2386_));
 sky130_fd_sc_hd__o32a_1 _6094_ (.A1(net174),
    .A2(_2385_),
    .A3(_2386_),
    .B1(_0789_),
    .B2(net88),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _6095_ (.A0(_2387_),
    .A1(net260),
    .S(net77),
    .X(_0276_));
 sky130_fd_sc_hd__nor2_1 _6096_ (.A(net166),
    .B(_0829_),
    .Y(_2388_));
 sky130_fd_sc_hd__a211o_1 _6097_ (.A1(net166),
    .A2(_0721_),
    .B1(_2325_),
    .C1(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__nor2_1 _6098_ (.A(net92),
    .B(_0829_),
    .Y(_2390_));
 sky130_fd_sc_hd__a211o_1 _6099_ (.A1(\as1802.regs[2][8] ),
    .A2(net92),
    .B1(_2390_),
    .C1(net94),
    .X(_2391_));
 sky130_fd_sc_hd__nand2_1 _6100_ (.A(_2389_),
    .B(_2391_),
    .Y(_2392_));
 sky130_fd_sc_hd__a221o_1 _6101_ (.A1(_3501_),
    .A2(_0720_),
    .B1(_2392_),
    .B2(_3528_),
    .C1(_2327_),
    .X(_2393_));
 sky130_fd_sc_hd__a21oi_1 _6102_ (.A1(_3623_),
    .A2(_2327_),
    .B1(net174),
    .Y(_2394_));
 sky130_fd_sc_hd__o2bb2a_1 _6103_ (.A1_N(_2393_),
    .A2_N(_2394_),
    .B1(_0721_),
    .B2(net88),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(_2395_),
    .A1(net292),
    .S(net77),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _6105_ (.A0(_0942_),
    .A1(_0963_),
    .S(net118),
    .X(_2396_));
 sky130_fd_sc_hd__inv_2 _6106_ (.A(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__nor2_1 _6107_ (.A(net93),
    .B(_0963_),
    .Y(_2398_));
 sky130_fd_sc_hd__a211o_1 _6108_ (.A1(\as1802.regs[2][9] ),
    .A2(net93),
    .B1(_2398_),
    .C1(net94),
    .X(_2399_));
 sky130_fd_sc_hd__o21a_1 _6109_ (.A1(_2325_),
    .A2(_2397_),
    .B1(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__o221a_1 _6110_ (.A1(net95),
    .A2(_0943_),
    .B1(_2400_),
    .B2(net96),
    .C1(net86),
    .X(_2401_));
 sky130_fd_sc_hd__nor2_1 _6111_ (.A(_3616_),
    .B(net86),
    .Y(_2402_));
 sky130_fd_sc_hd__o32a_1 _6112_ (.A1(net174),
    .A2(_2401_),
    .A3(_2402_),
    .B1(_0943_),
    .B2(net88),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _6113_ (.A0(_2403_),
    .A1(net290),
    .S(net77),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _6114_ (.A0(_0991_),
    .A1(_1011_),
    .S(net118),
    .X(_2404_));
 sky130_fd_sc_hd__inv_2 _6115_ (.A(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__nor2_1 _6116_ (.A(net92),
    .B(_1011_),
    .Y(_2406_));
 sky130_fd_sc_hd__a211o_1 _6117_ (.A1(\as1802.regs[2][10] ),
    .A2(net92),
    .B1(_2406_),
    .C1(net94),
    .X(_2407_));
 sky130_fd_sc_hd__o21a_1 _6118_ (.A1(_2325_),
    .A2(_2405_),
    .B1(_2407_),
    .X(_2408_));
 sky130_fd_sc_hd__o221a_1 _6119_ (.A1(net95),
    .A2(_0992_),
    .B1(_2408_),
    .B2(net96),
    .C1(net86),
    .X(_2409_));
 sky130_fd_sc_hd__nor2_1 _6120_ (.A(_0462_),
    .B(net86),
    .Y(_2410_));
 sky130_fd_sc_hd__o32a_1 _6121_ (.A1(net174),
    .A2(_2409_),
    .A3(_2410_),
    .B1(_0992_),
    .B2(net88),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_1 _6122_ (.A0(_2411_),
    .A1(net302),
    .S(net77),
    .X(_0279_));
 sky130_fd_sc_hd__and2b_1 _6123_ (.A_N(net88),
    .B(_1041_),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(_1041_),
    .A1(_1061_),
    .S(net118),
    .X(_2413_));
 sky130_fd_sc_hd__inv_2 _6125_ (.A(_2413_),
    .Y(_2414_));
 sky130_fd_sc_hd__nor2_1 _6126_ (.A(net92),
    .B(_1061_),
    .Y(_2415_));
 sky130_fd_sc_hd__a211o_1 _6127_ (.A1(\as1802.regs[2][11] ),
    .A2(net92),
    .B1(_2415_),
    .C1(net94),
    .X(_2416_));
 sky130_fd_sc_hd__o21ai_2 _6128_ (.A1(_2325_),
    .A2(_2414_),
    .B1(_2416_),
    .Y(_2417_));
 sky130_fd_sc_hd__a221o_1 _6129_ (.A1(_3501_),
    .A2(_1041_),
    .B1(_2417_),
    .B2(_3528_),
    .C1(_2327_),
    .X(_2418_));
 sky130_fd_sc_hd__or2_1 _6130_ (.A(_0472_),
    .B(net86),
    .X(_2419_));
 sky130_fd_sc_hd__a311o_1 _6131_ (.A1(_3432_),
    .A2(_2418_),
    .A3(_2419_),
    .B1(net77),
    .C1(_2412_),
    .X(_2420_));
 sky130_fd_sc_hd__a21bo_1 _6132_ (.A1(net282),
    .A2(net77),
    .B1_N(_2420_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _6133_ (.A0(_1086_),
    .A1(_1106_),
    .S(net118),
    .X(_2421_));
 sky130_fd_sc_hd__inv_2 _6134_ (.A(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__nor2_1 _6135_ (.A(net92),
    .B(_1106_),
    .Y(_2423_));
 sky130_fd_sc_hd__a211o_1 _6136_ (.A1(\as1802.regs[2][12] ),
    .A2(net92),
    .B1(_2423_),
    .C1(net94),
    .X(_2424_));
 sky130_fd_sc_hd__o21a_1 _6137_ (.A1(_2325_),
    .A2(_2422_),
    .B1(_2424_),
    .X(_2425_));
 sky130_fd_sc_hd__o221a_1 _6138_ (.A1(_3500_),
    .A2(_1087_),
    .B1(_2425_),
    .B2(net96),
    .C1(net86),
    .X(_2426_));
 sky130_fd_sc_hd__nor2_1 _6139_ (.A(_3608_),
    .B(net86),
    .Y(_2427_));
 sky130_fd_sc_hd__o32a_1 _6140_ (.A1(net174),
    .A2(_2426_),
    .A3(_2427_),
    .B1(_1087_),
    .B2(net88),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _6141_ (.A0(_2428_),
    .A1(net298),
    .S(net77),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _6142_ (.A0(_1135_),
    .A1(_1157_),
    .S(net118),
    .X(_2429_));
 sky130_fd_sc_hd__inv_2 _6143_ (.A(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__nor2_1 _6144_ (.A(net92),
    .B(_1157_),
    .Y(_2431_));
 sky130_fd_sc_hd__a211o_1 _6145_ (.A1(\as1802.regs[2][13] ),
    .A2(net92),
    .B1(_2431_),
    .C1(_0527_),
    .X(_2432_));
 sky130_fd_sc_hd__o21a_1 _6146_ (.A1(_2325_),
    .A2(_2430_),
    .B1(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__o221a_1 _6147_ (.A1(_3500_),
    .A2(_1136_),
    .B1(_2433_),
    .B2(net96),
    .C1(net86),
    .X(_2434_));
 sky130_fd_sc_hd__nor2_1 _6148_ (.A(_3600_),
    .B(net86),
    .Y(_2435_));
 sky130_fd_sc_hd__o32a_1 _6149_ (.A1(net174),
    .A2(_2434_),
    .A3(_2435_),
    .B1(_1136_),
    .B2(net88),
    .X(_2436_));
 sky130_fd_sc_hd__mux2_1 _6150_ (.A0(_2436_),
    .A1(net286),
    .S(net77),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _6151_ (.A0(_1183_),
    .A1(_1206_),
    .S(_3443_),
    .X(_2437_));
 sky130_fd_sc_hd__inv_2 _6152_ (.A(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__nor2_1 _6153_ (.A(net92),
    .B(_1206_),
    .Y(_2439_));
 sky130_fd_sc_hd__a211o_1 _6154_ (.A1(\as1802.regs[2][14] ),
    .A2(net92),
    .B1(_2439_),
    .C1(_0527_),
    .X(_2440_));
 sky130_fd_sc_hd__o21a_1 _6155_ (.A1(_2325_),
    .A2(_2438_),
    .B1(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__o221a_1 _6156_ (.A1(_3500_),
    .A2(_1184_),
    .B1(_2441_),
    .B2(_3527_),
    .C1(net86),
    .X(_2442_));
 sky130_fd_sc_hd__nor2_1 _6157_ (.A(_3592_),
    .B(net86),
    .Y(_2443_));
 sky130_fd_sc_hd__o32a_1 _6158_ (.A1(net174),
    .A2(_2442_),
    .A3(_2443_),
    .B1(_1184_),
    .B2(net88),
    .X(_2444_));
 sky130_fd_sc_hd__mux2_1 _6159_ (.A0(_2444_),
    .A1(net280),
    .S(net77),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _6160_ (.A0(_1227_),
    .A1(_1246_),
    .S(_3443_),
    .X(_2445_));
 sky130_fd_sc_hd__inv_2 _6161_ (.A(_2445_),
    .Y(_2446_));
 sky130_fd_sc_hd__nor2_1 _6162_ (.A(net93),
    .B(_1246_),
    .Y(_2447_));
 sky130_fd_sc_hd__a211o_1 _6163_ (.A1(\as1802.regs[2][15] ),
    .A2(net93),
    .B1(_2447_),
    .C1(_0527_),
    .X(_2448_));
 sky130_fd_sc_hd__o21a_1 _6164_ (.A1(_2325_),
    .A2(_2446_),
    .B1(_2448_),
    .X(_2449_));
 sky130_fd_sc_hd__o221a_1 _6165_ (.A1(_3500_),
    .A2(_1228_),
    .B1(_2449_),
    .B2(_3527_),
    .C1(net86),
    .X(_2450_));
 sky130_fd_sc_hd__nor2_1 _6166_ (.A(_0485_),
    .B(net87),
    .Y(_2451_));
 sky130_fd_sc_hd__o32a_1 _6167_ (.A1(net174),
    .A2(_2450_),
    .A3(_2451_),
    .B1(_1228_),
    .B2(net88),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _6168_ (.A0(_2452_),
    .A1(net306),
    .S(net77),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _6169_ (.A0(net292),
    .A1(net272),
    .S(_2310_),
    .X(_2453_));
 sky130_fd_sc_hd__or2_1 _6170_ (.A(net398),
    .B(_3547_),
    .X(_2454_));
 sky130_fd_sc_hd__o211a_1 _6171_ (.A1(_3548_),
    .A2(_2453_),
    .B1(_2454_),
    .C1(net212),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _6172_ (.A0(net290),
    .A1(net268),
    .S(_2310_),
    .X(_2455_));
 sky130_fd_sc_hd__or2_1 _6173_ (.A(net392),
    .B(_3547_),
    .X(_2456_));
 sky130_fd_sc_hd__o211a_1 _6174_ (.A1(_3548_),
    .A2(_2455_),
    .B1(_2456_),
    .C1(net212),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _6175_ (.A0(net302),
    .A1(net266),
    .S(_2310_),
    .X(_2457_));
 sky130_fd_sc_hd__or2_1 _6176_ (.A(net379),
    .B(_3547_),
    .X(_2458_));
 sky130_fd_sc_hd__o211a_1 _6177_ (.A1(_3548_),
    .A2(_2457_),
    .B1(_2458_),
    .C1(net212),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _6178_ (.A0(net282),
    .A1(net264),
    .S(_2310_),
    .X(_2459_));
 sky130_fd_sc_hd__or2_1 _6179_ (.A(net364),
    .B(_3547_),
    .X(_2460_));
 sky130_fd_sc_hd__o211a_1 _6180_ (.A1(_3548_),
    .A2(_2459_),
    .B1(_2460_),
    .C1(net212),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _6181_ (.A0(net298),
    .A1(net262),
    .S(_2310_),
    .X(_2461_));
 sky130_fd_sc_hd__or2_1 _6182_ (.A(net718),
    .B(_3547_),
    .X(_2462_));
 sky130_fd_sc_hd__o211a_1 _6183_ (.A1(_3548_),
    .A2(_2461_),
    .B1(_2462_),
    .C1(net212),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _6184_ (.A0(net286),
    .A1(net256),
    .S(_2310_),
    .X(_2463_));
 sky130_fd_sc_hd__or2_1 _6185_ (.A(net335),
    .B(_3547_),
    .X(_2464_));
 sky130_fd_sc_hd__o211a_1 _6186_ (.A1(_3548_),
    .A2(_2463_),
    .B1(net336),
    .C1(net212),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _6187_ (.A0(net280),
    .A1(net258),
    .S(_2310_),
    .X(_2465_));
 sky130_fd_sc_hd__or2_1 _6188_ (.A(net362),
    .B(_3547_),
    .X(_2466_));
 sky130_fd_sc_hd__o211a_1 _6189_ (.A1(_3548_),
    .A2(_2465_),
    .B1(_2466_),
    .C1(net212),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _6190_ (.A0(net306),
    .A1(net260),
    .S(_2310_),
    .X(_2467_));
 sky130_fd_sc_hd__or2_1 _6191_ (.A(net385),
    .B(_3547_),
    .X(_2468_));
 sky130_fd_sc_hd__o211a_1 _6192_ (.A1(_3548_),
    .A2(_2467_),
    .B1(_2468_),
    .C1(net212),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _6193_ (.A0(net333),
    .A1(net292),
    .S(_3550_),
    .X(_2469_));
 sky130_fd_sc_hd__or2_1 _6194_ (.A(_3464_),
    .B(net334),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(_3454_),
    .A1(_3455_),
    .S(_3550_),
    .X(_2470_));
 sky130_fd_sc_hd__nand2_1 _6196_ (.A(net212),
    .B(net372),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(_3452_),
    .A1(_3453_),
    .S(_3550_),
    .X(_2471_));
 sky130_fd_sc_hd__nand2_1 _6198_ (.A(net212),
    .B(net462),
    .Y(_0299_));
 sky130_fd_sc_hd__mux2_1 _6199_ (.A0(_3450_),
    .A1(_3451_),
    .S(_3550_),
    .X(_2472_));
 sky130_fd_sc_hd__nand2_1 _6200_ (.A(net213),
    .B(net374),
    .Y(_0300_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(_3448_),
    .A1(_3449_),
    .S(_3550_),
    .X(_2473_));
 sky130_fd_sc_hd__nand2_1 _6202_ (.A(net213),
    .B(net370),
    .Y(_0301_));
 sky130_fd_sc_hd__mux2_1 _6203_ (.A0(net340),
    .A1(net286),
    .S(_3550_),
    .X(_2474_));
 sky130_fd_sc_hd__or2_1 _6204_ (.A(_3464_),
    .B(net341),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _6205_ (.A0(net331),
    .A1(net280),
    .S(_3550_),
    .X(_2475_));
 sky130_fd_sc_hd__or2_1 _6206_ (.A(net206),
    .B(net332),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _6207_ (.A0(_3446_),
    .A1(_3447_),
    .S(_3550_),
    .X(_2476_));
 sky130_fd_sc_hd__nand2_1 _6208_ (.A(net213),
    .B(net378),
    .Y(_0304_));
 sky130_fd_sc_hd__a31o_1 _6209_ (.A1(net173),
    .A2(net104),
    .A3(_3535_),
    .B1(net830),
    .X(_2477_));
 sky130_fd_sc_hd__and3b_1 _6210_ (.A_N(_1255_),
    .B(net831),
    .C(net210),
    .X(_0305_));
 sky130_fd_sc_hd__nor2_1 _6211_ (.A(net45),
    .B(_3556_),
    .Y(_2478_));
 sky130_fd_sc_hd__a31o_1 _6212_ (.A1(net356),
    .A2(\as1802.mem_write ),
    .A3(_3481_),
    .B1(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__nand2_1 _6213_ (.A(net210),
    .B(net357),
    .Y(_0306_));
 sky130_fd_sc_hd__nand2_1 _6214_ (.A(net210),
    .B(_3544_),
    .Y(_2480_));
 sky130_fd_sc_hd__a21o_1 _6215_ (.A1(net270),
    .A2(_3543_),
    .B1(_2480_),
    .X(_0307_));
 sky130_fd_sc_hd__or3_1 _6216_ (.A(net356),
    .B(_3457_),
    .C(net352),
    .X(_2481_));
 sky130_fd_sc_hd__a22o_1 _6217_ (.A1(_3550_),
    .A2(_2307_),
    .B1(_2481_),
    .B2(net854),
    .X(_2482_));
 sky130_fd_sc_hd__and2_1 _6218_ (.A(net213),
    .B(_2482_),
    .X(_0308_));
 sky130_fd_sc_hd__a211o_1 _6219_ (.A1(net161),
    .A2(net315),
    .B1(_0514_),
    .C1(net117),
    .X(_2483_));
 sky130_fd_sc_hd__or4_1 _6220_ (.A(_3532_),
    .B(_3553_),
    .C(_0513_),
    .D(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__o21ai_1 _6221_ (.A1(_3570_),
    .A2(_2484_),
    .B1(net209),
    .Y(_2485_));
 sky130_fd_sc_hd__a21oi_1 _6222_ (.A1(_3445_),
    .A2(_2484_),
    .B1(_2485_),
    .Y(_0309_));
 sky130_fd_sc_hd__nand2_1 _6223_ (.A(_3442_),
    .B(_1567_),
    .Y(_2486_));
 sky130_fd_sc_hd__o211a_1 _6224_ (.A1(net35),
    .A2(_1567_),
    .B1(_2486_),
    .C1(net207),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _6225_ (.A(_3441_),
    .B(_1567_),
    .Y(_2487_));
 sky130_fd_sc_hd__o211a_1 _6226_ (.A1(net36),
    .A2(_1567_),
    .B1(_2487_),
    .C1(net209),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _6227_ (.A0(net809),
    .A1(net37),
    .S(_1566_),
    .X(_2488_));
 sky130_fd_sc_hd__or2_1 _6228_ (.A(net206),
    .B(_2488_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _6229_ (.A0(net827),
    .A1(net38),
    .S(_1566_),
    .X(_2489_));
 sky130_fd_sc_hd__or2_1 _6230_ (.A(net206),
    .B(_2489_),
    .X(_0317_));
 sky130_fd_sc_hd__o2bb2a_1 _6231_ (.A1_N(net865),
    .A2_N(_2292_),
    .B1(_2291_),
    .B2(_3553_),
    .X(_2490_));
 sky130_fd_sc_hd__nor2_1 _6232_ (.A(net206),
    .B(net866),
    .Y(_0318_));
 sky130_fd_sc_hd__nor2_1 _6233_ (.A(_3433_),
    .B(net139),
    .Y(_2491_));
 sky130_fd_sc_hd__nor2_1 _6234_ (.A(net120),
    .B(net139),
    .Y(_2492_));
 sky130_fd_sc_hd__or2_1 _6235_ (.A(net120),
    .B(net139),
    .X(_2493_));
 sky130_fd_sc_hd__nand2_4 _6236_ (.A(_2262_),
    .B(_2493_),
    .Y(_2494_));
 sky130_fd_sc_hd__inv_2 _6237_ (.A(_2494_),
    .Y(_2495_));
 sky130_fd_sc_hd__and2_1 _6238_ (.A(net123),
    .B(_3477_),
    .X(_2496_));
 sky130_fd_sc_hd__or2_2 _6239_ (.A(net123),
    .B(_3477_),
    .X(_2497_));
 sky130_fd_sc_hd__and2_1 _6240_ (.A(net126),
    .B(_3476_),
    .X(_2498_));
 sky130_fd_sc_hd__nor2_1 _6241_ (.A(net124),
    .B(_3476_),
    .Y(_2499_));
 sky130_fd_sc_hd__or2_1 _6242_ (.A(net126),
    .B(_3476_),
    .X(_2500_));
 sky130_fd_sc_hd__nand2_1 _6243_ (.A(net127),
    .B(_3475_),
    .Y(_2501_));
 sky130_fd_sc_hd__nor2_1 _6244_ (.A(net127),
    .B(_3475_),
    .Y(_2502_));
 sky130_fd_sc_hd__nand2_1 _6245_ (.A(_3434_),
    .B(net148),
    .Y(_2503_));
 sky130_fd_sc_hd__and2_2 _6246_ (.A(_2501_),
    .B(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__nand2_1 _6247_ (.A(_2501_),
    .B(_2503_),
    .Y(_2505_));
 sky130_fd_sc_hd__nand2_2 _6248_ (.A(net130),
    .B(net106),
    .Y(_2506_));
 sky130_fd_sc_hd__inv_2 _6249_ (.A(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__nor2_2 _6250_ (.A(net130),
    .B(net106),
    .Y(_2508_));
 sky130_fd_sc_hd__nor2_2 _6251_ (.A(_3436_),
    .B(net154),
    .Y(_2509_));
 sky130_fd_sc_hd__nor2_1 _6252_ (.A(net132),
    .B(net107),
    .Y(_2510_));
 sky130_fd_sc_hd__nand2_1 _6253_ (.A(_3436_),
    .B(net154),
    .Y(_2511_));
 sky130_fd_sc_hd__nor2_2 _6254_ (.A(_2509_),
    .B(_2510_),
    .Y(_2512_));
 sky130_fd_sc_hd__or2_2 _6255_ (.A(_2509_),
    .B(_2510_),
    .X(_2513_));
 sky130_fd_sc_hd__nand2_2 _6256_ (.A(net133),
    .B(net108),
    .Y(_2514_));
 sky130_fd_sc_hd__nor2_1 _6257_ (.A(net133),
    .B(net108),
    .Y(_2515_));
 sky130_fd_sc_hd__inv_2 _6258_ (.A(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__nand2_2 _6259_ (.A(_2514_),
    .B(_2516_),
    .Y(_2517_));
 sky130_fd_sc_hd__nor2_1 _6260_ (.A(net135),
    .B(net111),
    .Y(_2518_));
 sky130_fd_sc_hd__nand2_2 _6261_ (.A(_3438_),
    .B(net160),
    .Y(_2519_));
 sky130_fd_sc_hd__or2_2 _6262_ (.A(_2517_),
    .B(_2518_),
    .X(_2520_));
 sky130_fd_sc_hd__a21oi_1 _6263_ (.A1(_2514_),
    .A2(_2520_),
    .B1(_2513_),
    .Y(_2521_));
 sky130_fd_sc_hd__or2_1 _6264_ (.A(_2509_),
    .B(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__nand2b_1 _6265_ (.A_N(_2508_),
    .B(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__a21o_1 _6266_ (.A1(_2506_),
    .A2(_2523_),
    .B1(_2505_),
    .X(_2524_));
 sky130_fd_sc_hd__nand2_1 _6267_ (.A(_2501_),
    .B(_2524_),
    .Y(_2525_));
 sky130_fd_sc_hd__a21o_1 _6268_ (.A1(_2500_),
    .A2(_2525_),
    .B1(_2498_),
    .X(_2526_));
 sky130_fd_sc_hd__a21o_1 _6269_ (.A1(_2497_),
    .A2(_2526_),
    .B1(_2496_),
    .X(_2527_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(_2494_),
    .B(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__a21o_1 _6271_ (.A1(_2494_),
    .A2(_2527_),
    .B1(_2491_),
    .X(_2529_));
 sky130_fd_sc_hd__nor2_1 _6272_ (.A(net126),
    .B(net238),
    .Y(_2530_));
 sky130_fd_sc_hd__or2_1 _6273_ (.A(net124),
    .B(net145),
    .X(_2531_));
 sky130_fd_sc_hd__and2_2 _6274_ (.A(_2166_),
    .B(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__nand2_2 _6275_ (.A(_2166_),
    .B(_2531_),
    .Y(_2533_));
 sky130_fd_sc_hd__and2b_2 _6276_ (.A_N(_2496_),
    .B(_2497_),
    .X(_2534_));
 sky130_fd_sc_hd__inv_2 _6277_ (.A(_2534_),
    .Y(_2535_));
 sky130_fd_sc_hd__nand2_2 _6278_ (.A(net135),
    .B(net111),
    .Y(_2536_));
 sky130_fd_sc_hd__nor2_4 _6279_ (.A(_2507_),
    .B(_2508_),
    .Y(_2537_));
 sky130_fd_sc_hd__inv_2 _6280_ (.A(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__or4_1 _6281_ (.A(_2505_),
    .B(_2513_),
    .C(_2532_),
    .D(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__or4b_1 _6282_ (.A(_2495_),
    .B(_2535_),
    .C(_2539_),
    .D_N(_2536_),
    .X(_2540_));
 sky130_fd_sc_hd__o21ai_1 _6283_ (.A1(_2520_),
    .A2(_2540_),
    .B1(_2529_),
    .Y(_2541_));
 sky130_fd_sc_hd__a22o_1 _6284_ (.A1(_3513_),
    .A2(_2529_),
    .B1(_2541_),
    .B2(net97),
    .X(_2542_));
 sky130_fd_sc_hd__and2_1 _6285_ (.A(_2519_),
    .B(_2536_),
    .X(_2543_));
 sky130_fd_sc_hd__nand2_1 _6286_ (.A(_2519_),
    .B(_2536_),
    .Y(_2544_));
 sky130_fd_sc_hd__nand2_1 _6287_ (.A(net63),
    .B(_2543_),
    .Y(_2545_));
 sky130_fd_sc_hd__a21o_1 _6288_ (.A1(_2536_),
    .A2(_2545_),
    .B1(net157),
    .X(_2546_));
 sky130_fd_sc_hd__nand3_1 _6289_ (.A(net157),
    .B(_2536_),
    .C(_2545_),
    .Y(_2547_));
 sky130_fd_sc_hd__and3_1 _6290_ (.A(net133),
    .B(_2546_),
    .C(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a21boi_2 _6291_ (.A1(net133),
    .A2(_2547_),
    .B1_N(_2546_),
    .Y(_2549_));
 sky130_fd_sc_hd__o21ba_1 _6292_ (.A1(_2510_),
    .A2(_2549_),
    .B1_N(_2509_),
    .X(_2550_));
 sky130_fd_sc_hd__a21o_1 _6293_ (.A1(_2506_),
    .A2(_2550_),
    .B1(_2508_),
    .X(_2551_));
 sky130_fd_sc_hd__or2_1 _6294_ (.A(_2505_),
    .B(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__nand2_1 _6295_ (.A(_2501_),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__o21a_1 _6296_ (.A1(_2498_),
    .A2(_2553_),
    .B1(_2500_),
    .X(_2554_));
 sky130_fd_sc_hd__a21o_1 _6297_ (.A1(_2534_),
    .A2(_2554_),
    .B1(_2496_),
    .X(_2555_));
 sky130_fd_sc_hd__nand2_1 _6298_ (.A(_3433_),
    .B(net139),
    .Y(_2556_));
 sky130_fd_sc_hd__a2111oi_1 _6299_ (.A1(_2555_),
    .A2(_2556_),
    .B1(\as1802.cond_inv ),
    .C1(_3514_),
    .D1(_2491_),
    .Y(_2557_));
 sky130_fd_sc_hd__nand2_2 _6300_ (.A(net135),
    .B(net160),
    .Y(_2558_));
 sky130_fd_sc_hd__nand2_1 _6301_ (.A(net871),
    .B(_2544_),
    .Y(_2559_));
 sky130_fd_sc_hd__a21bo_1 _6302_ (.A1(_2558_),
    .A2(_2559_),
    .B1_N(_2517_),
    .X(_2560_));
 sky130_fd_sc_hd__a21o_1 _6303_ (.A1(_2092_),
    .A2(_2560_),
    .B1(_2512_),
    .X(_2561_));
 sky130_fd_sc_hd__a21o_1 _6304_ (.A1(_2036_),
    .A2(_2561_),
    .B1(_2537_),
    .X(_2562_));
 sky130_fd_sc_hd__a21oi_1 _6305_ (.A1(_1947_),
    .A2(_2562_),
    .B1(_2504_),
    .Y(_2563_));
 sky130_fd_sc_hd__nor2_1 _6306_ (.A(_2005_),
    .B(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__or2_1 _6307_ (.A(_2530_),
    .B(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__a21oi_1 _6308_ (.A1(_2166_),
    .A2(_2565_),
    .B1(_2534_),
    .Y(_2566_));
 sky130_fd_sc_hd__nor2_1 _6309_ (.A(_2221_),
    .B(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__a21oi_1 _6310_ (.A1(_2262_),
    .A2(_2567_),
    .B1(_2492_),
    .Y(_2568_));
 sky130_fd_sc_hd__or2_1 _6311_ (.A(net135),
    .B(net164),
    .X(_2569_));
 sky130_fd_sc_hd__o211a_1 _6312_ (.A1(net120),
    .A2(net117),
    .B1(_3517_),
    .C1(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__o31a_1 _6313_ (.A1(\as1802.cond_inv ),
    .A2(net170),
    .A3(_3444_),
    .B1(net168),
    .X(_2571_));
 sky130_fd_sc_hd__or3b_1 _6314_ (.A(_2557_),
    .B(_2570_),
    .C_N(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__a221o_1 _6315_ (.A1(net164),
    .A2(_2542_),
    .B1(_2568_),
    .B2(net101),
    .C1(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__nand2_1 _6316_ (.A(_2519_),
    .B(_2545_),
    .Y(_2574_));
 sky130_fd_sc_hd__a21o_1 _6317_ (.A1(_2514_),
    .A2(_2574_),
    .B1(_2515_),
    .X(_2575_));
 sky130_fd_sc_hd__and2b_1 _6318_ (.A_N(_2509_),
    .B(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__or2_1 _6319_ (.A(_2510_),
    .B(_2576_),
    .X(_2577_));
 sky130_fd_sc_hd__a21o_1 _6320_ (.A1(_2506_),
    .A2(_2577_),
    .B1(_2508_),
    .X(_2578_));
 sky130_fd_sc_hd__o211a_1 _6321_ (.A1(_2502_),
    .A2(_2578_),
    .B1(_2533_),
    .C1(_2501_),
    .X(_2579_));
 sky130_fd_sc_hd__nor2_1 _6322_ (.A(_2499_),
    .B(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__o21a_1 _6323_ (.A1(_2496_),
    .A2(_2580_),
    .B1(_2497_),
    .X(_2581_));
 sky130_fd_sc_hd__and2_1 _6324_ (.A(_2494_),
    .B(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__o311a_1 _6325_ (.A1(_2491_),
    .A2(_2571_),
    .A3(_2582_),
    .B1(_2573_),
    .C1(net100),
    .X(_2583_));
 sky130_fd_sc_hd__or4_1 _6326_ (.A(net119),
    .B(net169),
    .C(net100),
    .D(_0580_),
    .X(_2584_));
 sky130_fd_sc_hd__a21oi_1 _6327_ (.A1(net168),
    .A2(_2584_),
    .B1(_0524_),
    .Y(_2585_));
 sky130_fd_sc_hd__nand2_1 _6328_ (.A(net95),
    .B(_0525_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_1 _6329_ (.A(net99),
    .B(_2118_),
    .Y(_2587_));
 sky130_fd_sc_hd__o211ai_1 _6330_ (.A1(net167),
    .A2(net94),
    .B1(_0593_),
    .C1(_3432_),
    .Y(_2588_));
 sky130_fd_sc_hd__or4_1 _6331_ (.A(_0517_),
    .B(_0558_),
    .C(_2586_),
    .D(_2587_),
    .X(_2589_));
 sky130_fd_sc_hd__or3_1 _6332_ (.A(_2585_),
    .B(_2588_),
    .C(_2589_),
    .X(_2590_));
 sky130_fd_sc_hd__or3_1 _6333_ (.A(_3518_),
    .B(_2542_),
    .C(_2570_),
    .X(_2591_));
 sky130_fd_sc_hd__a21o_1 _6334_ (.A1(_2514_),
    .A2(_2516_),
    .B1(_2558_),
    .X(_2592_));
 sky130_fd_sc_hd__a21o_1 _6335_ (.A1(_2092_),
    .A2(_2592_),
    .B1(_2512_),
    .X(_2593_));
 sky130_fd_sc_hd__a21o_1 _6336_ (.A1(_2036_),
    .A2(_2593_),
    .B1(_2537_),
    .X(_2594_));
 sky130_fd_sc_hd__a21oi_1 _6337_ (.A1(_1947_),
    .A2(_2594_),
    .B1(_2504_),
    .Y(_2595_));
 sky130_fd_sc_hd__nor2_1 _6338_ (.A(_2005_),
    .B(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__or2_1 _6339_ (.A(_2530_),
    .B(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__a21oi_1 _6340_ (.A1(_2166_),
    .A2(_2597_),
    .B1(_2534_),
    .Y(_2598_));
 sky130_fd_sc_hd__nor2_1 _6341_ (.A(_2221_),
    .B(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__o211ai_1 _6342_ (.A1(_2492_),
    .A2(_2599_),
    .B1(_3518_),
    .C1(_2262_),
    .Y(_2600_));
 sky130_fd_sc_hd__a31o_1 _6343_ (.A1(_0513_),
    .A2(_2591_),
    .A3(_2600_),
    .B1(_2583_),
    .X(_2601_));
 sky130_fd_sc_hd__mux2_1 _6344_ (.A0(_2601_),
    .A1(net871),
    .S(_2590_),
    .X(_2602_));
 sky130_fd_sc_hd__and2_1 _6345_ (.A(net210),
    .B(_2602_),
    .X(_0319_));
 sky130_fd_sc_hd__a32o_1 _6346_ (.A1(net105),
    .A2(_3579_),
    .A3(_0678_),
    .B1(_3553_),
    .B2(net161),
    .X(_2603_));
 sky130_fd_sc_hd__and2_1 _6347_ (.A(net207),
    .B(_2603_),
    .X(_0320_));
 sky130_fd_sc_hd__a41o_1 _6348_ (.A1(_3432_),
    .A2(_3440_),
    .A3(_3441_),
    .A4(net163),
    .B1(net102),
    .X(_2604_));
 sky130_fd_sc_hd__nor2_1 _6349_ (.A(_2318_),
    .B(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__o21ai_1 _6350_ (.A1(_0587_),
    .A2(_2283_),
    .B1(_3540_),
    .Y(_2606_));
 sky130_fd_sc_hd__nand2_1 _6351_ (.A(_2605_),
    .B(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__a21o_1 _6352_ (.A1(net833),
    .A2(_2607_),
    .B1(net206),
    .X(_2608_));
 sky130_fd_sc_hd__a41o_1 _6353_ (.A1(_3432_),
    .A2(_3576_),
    .A3(_2605_),
    .A4(_2606_),
    .B1(net834),
    .X(_0321_));
 sky130_fd_sc_hd__nor2_1 _6354_ (.A(net164),
    .B(_0500_),
    .Y(_2609_));
 sky130_fd_sc_hd__o21a_1 _6355_ (.A1(_2283_),
    .A2(_2609_),
    .B1(_3540_),
    .X(_2610_));
 sky130_fd_sc_hd__nor2_1 _6356_ (.A(net172),
    .B(net91),
    .Y(_2611_));
 sky130_fd_sc_hd__or4b_4 _6357_ (.A(_3541_),
    .B(_2610_),
    .C(_2611_),
    .D_N(_2605_),
    .X(_2612_));
 sky130_fd_sc_hd__mux2_1 _6358_ (.A0(net284),
    .A1(net354),
    .S(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__and2_1 _6359_ (.A(net207),
    .B(net355),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _6360_ (.A0(\as1802.P[1] ),
    .A1(net346),
    .S(_2612_),
    .X(_2614_));
 sky130_fd_sc_hd__and2_1 _6361_ (.A(net207),
    .B(net347),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _6362_ (.A0(\as1802.P[2] ),
    .A1(net350),
    .S(_2612_),
    .X(_2615_));
 sky130_fd_sc_hd__and2_1 _6363_ (.A(net207),
    .B(net351),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _6364_ (.A0(net310),
    .A1(net342),
    .S(_2612_),
    .X(_2616_));
 sky130_fd_sc_hd__and2_1 _6365_ (.A(net207),
    .B(net343),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _6366_ (.A0(\as1802.X[0] ),
    .A1(net344),
    .S(_2612_),
    .X(_2617_));
 sky130_fd_sc_hd__and2_1 _6367_ (.A(net207),
    .B(net345),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _6368_ (.A0(net278),
    .A1(net360),
    .S(_2612_),
    .X(_2618_));
 sky130_fd_sc_hd__and2_1 _6369_ (.A(net207),
    .B(net361),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _6370_ (.A0(\as1802.X[2] ),
    .A1(net358),
    .S(_2612_),
    .X(_2619_));
 sky130_fd_sc_hd__and2_1 _6371_ (.A(net207),
    .B(net359),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _6372_ (.A0(\as1802.X[3] ),
    .A1(net348),
    .S(_2612_),
    .X(_2620_));
 sky130_fd_sc_hd__and2_1 _6373_ (.A(net207),
    .B(net349),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _6374_ (.A(_3432_),
    .B(_0538_),
    .Y(_2621_));
 sky130_fd_sc_hd__or4b_1 _6375_ (.A(net96),
    .B(_2621_),
    .C(_0516_),
    .D_N(_0540_),
    .X(_2622_));
 sky130_fd_sc_hd__a2111o_2 _6376_ (.A1(net104),
    .A2(_2622_),
    .B1(_1566_),
    .C1(_3550_),
    .D1(_3549_),
    .X(_2623_));
 sky130_fd_sc_hd__a21o_1 _6377_ (.A1(_3511_),
    .A2(_3561_),
    .B1(_3577_),
    .X(_2624_));
 sky130_fd_sc_hd__o21ai_1 _6378_ (.A1(_2283_),
    .A2(_2624_),
    .B1(_0590_),
    .Y(_2625_));
 sky130_fd_sc_hd__a211o_1 _6379_ (.A1(net276),
    .A2(_3545_),
    .B1(_3558_),
    .C1(_0680_),
    .X(_2626_));
 sky130_fd_sc_hd__a31o_1 _6380_ (.A1(net164),
    .A2(net104),
    .A3(_0678_),
    .B1(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__a211o_4 _6381_ (.A1(_0541_),
    .A2(_2625_),
    .B1(_2627_),
    .C1(_2623_),
    .X(_2628_));
 sky130_fd_sc_hd__a22o_1 _6382_ (.A1(net354),
    .A2(_3579_),
    .B1(net91),
    .B2(net284),
    .X(_2629_));
 sky130_fd_sc_hd__nand2_2 _6383_ (.A(_3526_),
    .B(_3577_),
    .Y(_2630_));
 sky130_fd_sc_hd__a22o_1 _6384_ (.A1(_3526_),
    .A2(_2629_),
    .B1(_2630_),
    .B2(net135),
    .X(_2631_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(net31),
    .A1(_2631_),
    .S(net105),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _6386_ (.A0(_2632_),
    .A1(net855),
    .S(_2628_),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _6387_ (.A1(net346),
    .A2(_3579_),
    .B1(net91),
    .B2(net742),
    .X(_2633_));
 sky130_fd_sc_hd__a22o_1 _6388_ (.A1(net133),
    .A2(_2630_),
    .B1(_2633_),
    .B2(_3526_),
    .X(_2634_));
 sky130_fd_sc_hd__mux2_1 _6389_ (.A0(net32),
    .A1(_2634_),
    .S(net105),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_1 _6390_ (.A0(_2635_),
    .A1(net828),
    .S(_2628_),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _6391_ (.A1(net350),
    .A2(_3579_),
    .B1(net91),
    .B2(net776),
    .X(_2636_));
 sky130_fd_sc_hd__a22o_1 _6392_ (.A1(net132),
    .A2(_2630_),
    .B1(_2636_),
    .B2(_3526_),
    .X(_2637_));
 sky130_fd_sc_hd__mux2_1 _6393_ (.A0(net33),
    .A1(_2637_),
    .S(net105),
    .X(_2638_));
 sky130_fd_sc_hd__mux2_1 _6394_ (.A0(_2638_),
    .A1(net878),
    .S(_2628_),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _6395_ (.A1(net342),
    .A2(_3579_),
    .B1(net91),
    .B2(net310),
    .X(_2639_));
 sky130_fd_sc_hd__a22o_1 _6396_ (.A1(net130),
    .A2(_2630_),
    .B1(_2639_),
    .B2(_3526_),
    .X(_2640_));
 sky130_fd_sc_hd__mux2_1 _6397_ (.A0(net34),
    .A1(_2640_),
    .S(net105),
    .X(_2641_));
 sky130_fd_sc_hd__mux2_1 _6398_ (.A0(_2641_),
    .A1(net849),
    .S(_2628_),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _6399_ (.A1(net344),
    .A2(_3579_),
    .B1(net91),
    .B2(net431),
    .X(_2642_));
 sky130_fd_sc_hd__a22o_1 _6400_ (.A1(net127),
    .A2(_2630_),
    .B1(_2642_),
    .B2(_3526_),
    .X(_2643_));
 sky130_fd_sc_hd__mux2_1 _6401_ (.A0(net35),
    .A1(_2643_),
    .S(net105),
    .X(_2644_));
 sky130_fd_sc_hd__mux2_1 _6402_ (.A0(_2644_),
    .A1(net876),
    .S(_2628_),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _6403_ (.A1(net360),
    .A2(_3579_),
    .B1(net91),
    .B2(net278),
    .X(_2645_));
 sky130_fd_sc_hd__a22o_1 _6404_ (.A1(net126),
    .A2(_2630_),
    .B1(_2645_),
    .B2(_3526_),
    .X(_2646_));
 sky130_fd_sc_hd__mux2_1 _6405_ (.A0(net36),
    .A1(_2646_),
    .S(net105),
    .X(_2647_));
 sky130_fd_sc_hd__mux2_1 _6406_ (.A0(_2647_),
    .A1(net238),
    .S(_2628_),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _6407_ (.A1(net358),
    .A2(_3579_),
    .B1(net91),
    .B2(net819),
    .X(_2648_));
 sky130_fd_sc_hd__a22o_1 _6408_ (.A1(net123),
    .A2(_2630_),
    .B1(_2648_),
    .B2(_3526_),
    .X(_2649_));
 sky130_fd_sc_hd__mux2_1 _6409_ (.A0(net37),
    .A1(_2649_),
    .S(net105),
    .X(_2650_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(_2650_),
    .A1(net859),
    .S(_2628_),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _6411_ (.A1(net348),
    .A2(_3579_),
    .B1(net91),
    .B2(net472),
    .X(_2651_));
 sky130_fd_sc_hd__a22o_1 _6412_ (.A1(net120),
    .A2(_2630_),
    .B1(_2651_),
    .B2(_3526_),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_1 _6413_ (.A0(net38),
    .A1(_2652_),
    .S(net105),
    .X(_2653_));
 sky130_fd_sc_hd__mux2_1 _6414_ (.A0(_2653_),
    .A1(net533),
    .S(_2628_),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _6415_ (.A(_3579_),
    .B(_0678_),
    .Y(_2654_));
 sky130_fd_sc_hd__nand2_1 _6416_ (.A(_0590_),
    .B(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__or3b_1 _6417_ (.A(_3532_),
    .B(net172),
    .C_N(_3530_),
    .X(_2656_));
 sky130_fd_sc_hd__o21ai_1 _6418_ (.A1(net172),
    .A2(_3499_),
    .B1(_0679_),
    .Y(_2657_));
 sky130_fd_sc_hd__or4b_4 _6419_ (.A(_2604_),
    .B(_2655_),
    .C(_2657_),
    .D_N(_2656_),
    .X(_2658_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(net321),
    .B(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__or3_1 _6421_ (.A(net174),
    .B(_3444_),
    .C(_2658_),
    .X(_2660_));
 sky130_fd_sc_hd__a21oi_1 _6422_ (.A1(net322),
    .A2(_2660_),
    .B1(_3464_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(net324),
    .B(_2658_),
    .Y(_2661_));
 sky130_fd_sc_hd__or3b_1 _6424_ (.A(_2658_),
    .B(net174),
    .C_N(net169),
    .X(_2662_));
 sky130_fd_sc_hd__a21oi_1 _6425_ (.A1(net325),
    .A2(_2662_),
    .B1(_3464_),
    .Y(_0343_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(net312),
    .B(_2658_),
    .Y(_2663_));
 sky130_fd_sc_hd__or3b_1 _6427_ (.A(_2658_),
    .B(net174),
    .C_N(net168),
    .X(_2664_));
 sky130_fd_sc_hd__a21oi_1 _6428_ (.A1(net313),
    .A2(_2664_),
    .B1(_3464_),
    .Y(_0344_));
 sky130_fd_sc_hd__o21ai_1 _6429_ (.A1(_3442_),
    .A2(_3623_),
    .B1(_0535_),
    .Y(_2665_));
 sky130_fd_sc_hd__nand2_1 _6430_ (.A(_1931_),
    .B(_1935_),
    .Y(_2666_));
 sky130_fd_sc_hd__xor2_1 _6431_ (.A(_1876_),
    .B(_2666_),
    .X(_2667_));
 sky130_fd_sc_hd__mux2_1 _6432_ (.A0(_1875_),
    .A1(_2667_),
    .S(net228),
    .X(_2668_));
 sky130_fd_sc_hd__o221a_4 _6433_ (.A1(_1878_),
    .A2(net228),
    .B1(_2668_),
    .B2(net138),
    .C1(_1797_),
    .X(_2669_));
 sky130_fd_sc_hd__xnor2_1 _6434_ (.A(_3478_),
    .B(_2668_),
    .Y(_2670_));
 sky130_fd_sc_hd__inv_2 _6435_ (.A(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__o21a_1 _6436_ (.A1(_1887_),
    .A2(_1930_),
    .B1(_1886_),
    .X(_2672_));
 sky130_fd_sc_hd__nand2_1 _6437_ (.A(_1891_),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__o21a_1 _6438_ (.A1(_1891_),
    .A2(_2672_),
    .B1(_1938_),
    .X(_2674_));
 sky130_fd_sc_hd__o2bb2a_2 _6439_ (.A1_N(_2674_),
    .A2_N(_2673_),
    .B1(_1938_),
    .B2(_1890_),
    .X(_2675_));
 sky130_fd_sc_hd__nor2_1 _6440_ (.A(net141),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__inv_2 _6441_ (.A(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__xnor2_1 _6442_ (.A(_1887_),
    .B(_1930_),
    .Y(_2678_));
 sky130_fd_sc_hd__mux2_1 _6443_ (.A0(_1885_),
    .A1(_2678_),
    .S(_1938_),
    .X(_2679_));
 sky130_fd_sc_hd__nor2_1 _6444_ (.A(net244),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__nand2_1 _6445_ (.A(net250),
    .B(_2679_),
    .Y(_2681_));
 sky130_fd_sc_hd__nand2b_1 _6446_ (.A_N(_2680_),
    .B(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__o21ai_1 _6447_ (.A1(_1909_),
    .A2(_1921_),
    .B1(_1908_),
    .Y(_2683_));
 sky130_fd_sc_hd__xnor2_1 _6448_ (.A(_1925_),
    .B(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__mux2_2 _6449_ (.A0(_1899_),
    .A1(_2684_),
    .S(_1938_),
    .X(_2685_));
 sky130_fd_sc_hd__or2_1 _6450_ (.A(net146),
    .B(_2685_),
    .X(_2686_));
 sky130_fd_sc_hd__xnor2_1 _6451_ (.A(_1910_),
    .B(_1921_),
    .Y(_2687_));
 sky130_fd_sc_hd__mux2_1 _6452_ (.A0(_1906_),
    .A1(_2687_),
    .S(_1938_),
    .X(_2688_));
 sky130_fd_sc_hd__or2_1 _6453_ (.A(net150),
    .B(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__xnor2_2 _6454_ (.A(net150),
    .B(_2688_),
    .Y(_2690_));
 sky130_fd_sc_hd__a31o_1 _6455_ (.A1(_1932_),
    .A2(_1933_),
    .A3(_1937_),
    .B1(_1918_),
    .X(_2691_));
 sky130_fd_sc_hd__o211ai_2 _6456_ (.A1(_1882_),
    .A2(_1931_),
    .B1(_1937_),
    .C1(_3462_),
    .Y(_2692_));
 sky130_fd_sc_hd__and3_1 _6457_ (.A(net109),
    .B(_2691_),
    .C(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__a21oi_1 _6458_ (.A1(_2691_),
    .A2(_2692_),
    .B1(net109),
    .Y(_2694_));
 sky130_fd_sc_hd__or2_1 _6459_ (.A(_2693_),
    .B(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__nor2_1 _6460_ (.A(net121),
    .B(net110),
    .Y(_2696_));
 sky130_fd_sc_hd__or3_4 _6461_ (.A(_2693_),
    .B(_2694_),
    .C(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__xor2_1 _6462_ (.A(_1915_),
    .B(_1920_),
    .X(_2698_));
 sky130_fd_sc_hd__mux2_4 _6463_ (.A0(_1912_),
    .A1(_2698_),
    .S(_1938_),
    .X(_2699_));
 sky130_fd_sc_hd__nor2_1 _6464_ (.A(net153),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__o21ba_1 _6465_ (.A1(net153),
    .A2(_2699_),
    .B1_N(_2693_),
    .X(_2701_));
 sky130_fd_sc_hd__and2_1 _6466_ (.A(_2697_),
    .B(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__and2_1 _6467_ (.A(net153),
    .B(_2699_),
    .X(_2703_));
 sky130_fd_sc_hd__nor3_1 _6468_ (.A(_2690_),
    .B(_2702_),
    .C(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__o31a_1 _6469_ (.A1(_2690_),
    .A2(_2702_),
    .A3(_2703_),
    .B1(_2689_),
    .X(_2705_));
 sky130_fd_sc_hd__a21o_1 _6470_ (.A1(net146),
    .A2(_2685_),
    .B1(_2689_),
    .X(_2706_));
 sky130_fd_sc_hd__xnor2_1 _6471_ (.A(net146),
    .B(_2685_),
    .Y(_2707_));
 sky130_fd_sc_hd__a2111o_1 _6472_ (.A1(_2697_),
    .A2(_2701_),
    .B1(_2703_),
    .C1(_2707_),
    .D1(_2690_),
    .X(_2708_));
 sky130_fd_sc_hd__a31oi_1 _6473_ (.A1(_2686_),
    .A2(_2706_),
    .A3(_2708_),
    .B1(_2682_),
    .Y(_2709_));
 sky130_fd_sc_hd__or2_1 _6474_ (.A(_2680_),
    .B(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__a21bo_1 _6475_ (.A1(net141),
    .A2(_2675_),
    .B1_N(_2680_),
    .X(_2711_));
 sky130_fd_sc_hd__xnor2_1 _6476_ (.A(net141),
    .B(_2675_),
    .Y(_2712_));
 sky130_fd_sc_hd__a311o_1 _6477_ (.A1(_2686_),
    .A2(_2706_),
    .A3(_2708_),
    .B1(_2712_),
    .C1(_2682_),
    .X(_2713_));
 sky130_fd_sc_hd__a31o_4 _6478_ (.A1(_2677_),
    .A2(_2711_),
    .A3(_2713_),
    .B1(_2671_),
    .X(_2714_));
 sky130_fd_sc_hd__nand2_4 _6479_ (.A(_2669_),
    .B(net233),
    .Y(_2715_));
 sky130_fd_sc_hd__xor2_1 _6480_ (.A(_2710_),
    .B(_2712_),
    .X(_2716_));
 sky130_fd_sc_hd__mux2_1 _6481_ (.A0(_2675_),
    .A1(_2716_),
    .S(_2715_),
    .X(_2717_));
 sky130_fd_sc_hd__nor2_1 _6482_ (.A(net138),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__nand2_1 _6483_ (.A(net138),
    .B(_2717_),
    .Y(_2719_));
 sky130_fd_sc_hd__xnor2_1 _6484_ (.A(_3478_),
    .B(_2717_),
    .Y(_2720_));
 sky130_fd_sc_hd__and4_1 _6485_ (.A(_2682_),
    .B(_2686_),
    .C(_2706_),
    .D(_2708_),
    .X(_2721_));
 sky130_fd_sc_hd__or2_1 _6486_ (.A(_2709_),
    .B(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__and3_1 _6487_ (.A(_2669_),
    .B(_2679_),
    .C(net233),
    .X(_2723_));
 sky130_fd_sc_hd__a21oi_2 _6488_ (.A1(_2715_),
    .A2(_2722_),
    .B1(_2723_),
    .Y(_2724_));
 sky130_fd_sc_hd__inv_2 _6489_ (.A(_2724_),
    .Y(_2725_));
 sky130_fd_sc_hd__and2_1 _6490_ (.A(_3477_),
    .B(_2724_),
    .X(_2726_));
 sky130_fd_sc_hd__o21a_1 _6491_ (.A1(_2702_),
    .A2(_2703_),
    .B1(_2690_),
    .X(_2727_));
 sky130_fd_sc_hd__a211o_1 _6492_ (.A1(_2669_),
    .A2(_2714_),
    .B1(_2727_),
    .C1(_2704_),
    .X(_2728_));
 sky130_fd_sc_hd__nand3b_2 _6493_ (.A_N(_2688_),
    .B(_2714_),
    .C(_2669_),
    .Y(_2729_));
 sky130_fd_sc_hd__nand2_1 _6494_ (.A(_2728_),
    .B(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__a21oi_2 _6495_ (.A1(_2728_),
    .A2(_2729_),
    .B1(net146),
    .Y(_2731_));
 sky130_fd_sc_hd__and3_1 _6496_ (.A(net146),
    .B(_2728_),
    .C(_2729_),
    .X(_2732_));
 sky130_fd_sc_hd__nor2_1 _6497_ (.A(_2731_),
    .B(_2732_),
    .Y(_2733_));
 sky130_fd_sc_hd__xnor2_1 _6498_ (.A(_2705_),
    .B(_2707_),
    .Y(_2734_));
 sky130_fd_sc_hd__nand3b_1 _6499_ (.A_N(_2685_),
    .B(_2714_),
    .C(_2669_),
    .Y(_2735_));
 sky130_fd_sc_hd__a21o_1 _6500_ (.A1(_2669_),
    .A2(_2714_),
    .B1(_2734_),
    .X(_2736_));
 sky130_fd_sc_hd__and2_1 _6501_ (.A(_2735_),
    .B(_2736_),
    .X(_2737_));
 sky130_fd_sc_hd__a21oi_2 _6502_ (.A1(_2735_),
    .A2(_2736_),
    .B1(net244),
    .Y(_2738_));
 sky130_fd_sc_hd__and3_1 _6503_ (.A(net244),
    .B(_2735_),
    .C(_2736_),
    .X(_2739_));
 sky130_fd_sc_hd__nor2_1 _6504_ (.A(_2738_),
    .B(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__or4_4 _6505_ (.A(_2731_),
    .B(_2732_),
    .C(_2738_),
    .D(_2739_),
    .X(_2741_));
 sky130_fd_sc_hd__or2_1 _6506_ (.A(_2700_),
    .B(_2703_),
    .X(_2742_));
 sky130_fd_sc_hd__nand2b_1 _6507_ (.A_N(_2693_),
    .B(_2697_),
    .Y(_2743_));
 sky130_fd_sc_hd__xor2_1 _6508_ (.A(_2742_),
    .B(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__nand3b_1 _6509_ (.A_N(_2699_),
    .B(net233),
    .C(_2669_),
    .Y(_2745_));
 sky130_fd_sc_hd__a21o_1 _6510_ (.A1(_2669_),
    .A2(net233),
    .B1(_2744_),
    .X(_2746_));
 sky130_fd_sc_hd__and2_1 _6511_ (.A(_2745_),
    .B(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__a21oi_1 _6512_ (.A1(_2745_),
    .A2(_2746_),
    .B1(net150),
    .Y(_2748_));
 sky130_fd_sc_hd__nand3_1 _6513_ (.A(net150),
    .B(_2745_),
    .C(_2746_),
    .Y(_2749_));
 sky130_fd_sc_hd__nand2b_1 _6514_ (.A_N(_2748_),
    .B(_2749_),
    .Y(_2750_));
 sky130_fd_sc_hd__a21oi_1 _6515_ (.A1(_2669_),
    .A2(_2714_),
    .B1(net110),
    .Y(_2751_));
 sky130_fd_sc_hd__xnor2_2 _6516_ (.A(net121),
    .B(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__or2_1 _6517_ (.A(net155),
    .B(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__nand2_1 _6518_ (.A(net155),
    .B(_2752_),
    .Y(_2754_));
 sky130_fd_sc_hd__nor2_1 _6519_ (.A(net122),
    .B(net110),
    .Y(_2755_));
 sky130_fd_sc_hd__a21o_1 _6520_ (.A1(net155),
    .A2(_2752_),
    .B1(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__and4_1 _6521_ (.A(_2669_),
    .B(_2691_),
    .C(_2692_),
    .D(_2714_),
    .X(_2757_));
 sky130_fd_sc_hd__nand2_1 _6522_ (.A(_2695_),
    .B(_2696_),
    .Y(_2758_));
 sky130_fd_sc_hd__a31o_1 _6523_ (.A1(_2697_),
    .A2(_2715_),
    .A3(_2758_),
    .B1(_2757_),
    .X(_2759_));
 sky130_fd_sc_hd__xnor2_1 _6524_ (.A(net107),
    .B(_2759_),
    .Y(_2760_));
 sky130_fd_sc_hd__a21o_1 _6525_ (.A1(_2753_),
    .A2(_2756_),
    .B1(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__nor2_1 _6526_ (.A(_2750_),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__a2111o_1 _6527_ (.A1(_2753_),
    .A2(_2756_),
    .B1(_2760_),
    .C1(_2750_),
    .D1(_2741_),
    .X(_2763_));
 sky130_fd_sc_hd__a31o_1 _6528_ (.A1(net107),
    .A2(_2749_),
    .A3(_2759_),
    .B1(_2748_),
    .X(_2764_));
 sky130_fd_sc_hd__and2b_1 _6529_ (.A_N(_2739_),
    .B(_2731_),
    .X(_2765_));
 sky130_fd_sc_hd__a311oi_2 _6530_ (.A1(_2733_),
    .A2(_2740_),
    .A3(_2764_),
    .B1(_2765_),
    .C1(_2738_),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_1 _6531_ (.A(_2763_),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__xnor2_1 _6532_ (.A(net141),
    .B(_2724_),
    .Y(_2768_));
 sky130_fd_sc_hd__a21o_1 _6533_ (.A1(_2767_),
    .A2(_2768_),
    .B1(_2726_),
    .X(_2769_));
 sky130_fd_sc_hd__nor2_1 _6534_ (.A(_2720_),
    .B(_2769_),
    .Y(_2770_));
 sky130_fd_sc_hd__nand2_1 _6535_ (.A(_2720_),
    .B(_2768_),
    .Y(_2771_));
 sky130_fd_sc_hd__a21o_1 _6536_ (.A1(_2763_),
    .A2(_2766_),
    .B1(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__a21oi_1 _6537_ (.A1(_2719_),
    .A2(_2726_),
    .B1(_2718_),
    .Y(_2773_));
 sky130_fd_sc_hd__a41oi_1 _6538_ (.A1(_2671_),
    .A2(_2677_),
    .A3(_2711_),
    .A4(_2713_),
    .B1(_2669_),
    .Y(_2774_));
 sky130_fd_sc_hd__o2bb2a_1 _6539_ (.A1_N(_2774_),
    .A2_N(net233),
    .B1(_2668_),
    .B2(_2715_),
    .X(_2775_));
 sky130_fd_sc_hd__and3_1 _6540_ (.A(_1797_),
    .B(_2773_),
    .C(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__nand2_4 _6541_ (.A(_2772_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__a21bo_1 _6542_ (.A1(_2720_),
    .A2(_2769_),
    .B1_N(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__o22a_1 _6543_ (.A1(_2717_),
    .A2(_2777_),
    .B1(_2778_),
    .B2(_2770_),
    .X(_2779_));
 sky130_fd_sc_hd__inv_2 _6544_ (.A(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__xnor2_1 _6545_ (.A(_2767_),
    .B(_2768_),
    .Y(_2781_));
 sky130_fd_sc_hd__mux2_1 _6546_ (.A0(_2725_),
    .A1(_2781_),
    .S(_2777_),
    .X(_2782_));
 sky130_fd_sc_hd__or2_1 _6547_ (.A(net138),
    .B(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__inv_2 _6548_ (.A(_2783_),
    .Y(_2784_));
 sky130_fd_sc_hd__o21a_1 _6549_ (.A1(_2762_),
    .A2(_2764_),
    .B1(_2733_),
    .X(_2785_));
 sky130_fd_sc_hd__o21ai_1 _6550_ (.A1(_2731_),
    .A2(_2785_),
    .B1(_2740_),
    .Y(_2786_));
 sky130_fd_sc_hd__o31a_1 _6551_ (.A1(_2731_),
    .A2(_2740_),
    .A3(_2785_),
    .B1(_2777_),
    .X(_2787_));
 sky130_fd_sc_hd__a2bb2o_1 _6552_ (.A1_N(_2737_),
    .A2_N(_2777_),
    .B1(_2786_),
    .B2(_2787_),
    .X(_2788_));
 sky130_fd_sc_hd__inv_2 _6553_ (.A(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__nand2_1 _6554_ (.A(_3477_),
    .B(_2788_),
    .Y(_2790_));
 sky130_fd_sc_hd__inv_2 _6555_ (.A(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__or2_1 _6556_ (.A(_3477_),
    .B(_2788_),
    .X(_2792_));
 sky130_fd_sc_hd__nor3_1 _6557_ (.A(_2733_),
    .B(_2762_),
    .C(_2764_),
    .Y(_2793_));
 sky130_fd_sc_hd__nor2_1 _6558_ (.A(_2785_),
    .B(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__mux2_2 _6559_ (.A0(_2730_),
    .A1(_2794_),
    .S(_2777_),
    .X(_2795_));
 sky130_fd_sc_hd__and2_1 _6560_ (.A(_3476_),
    .B(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__xnor2_2 _6561_ (.A(net244),
    .B(_2795_),
    .Y(_2797_));
 sky130_fd_sc_hd__a21bo_1 _6562_ (.A1(net107),
    .A2(_2759_),
    .B1_N(_2761_),
    .X(_2798_));
 sky130_fd_sc_hd__xor2_1 _6563_ (.A(_2750_),
    .B(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__mux2_1 _6564_ (.A0(_2747_),
    .A1(_2799_),
    .S(_2777_),
    .X(_2800_));
 sky130_fd_sc_hd__inv_2 _6565_ (.A(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__or2_2 _6566_ (.A(net146),
    .B(_2800_),
    .X(_2802_));
 sky130_fd_sc_hd__inv_2 _6567_ (.A(_2802_),
    .Y(_2803_));
 sky130_fd_sc_hd__and2_1 _6568_ (.A(net146),
    .B(_2800_),
    .X(_2804_));
 sky130_fd_sc_hd__nand3_1 _6569_ (.A(_2753_),
    .B(_2756_),
    .C(_2760_),
    .Y(_2805_));
 sky130_fd_sc_hd__and2_1 _6570_ (.A(_2761_),
    .B(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__mux2_1 _6571_ (.A0(_2759_),
    .A1(_2806_),
    .S(_2777_),
    .X(_2807_));
 sky130_fd_sc_hd__and2_1 _6572_ (.A(net106),
    .B(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__xnor2_1 _6573_ (.A(net150),
    .B(_2807_),
    .Y(_2809_));
 sky130_fd_sc_hd__inv_2 _6574_ (.A(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__and2_1 _6575_ (.A(_2753_),
    .B(_2754_),
    .X(_2811_));
 sky130_fd_sc_hd__xor2_1 _6576_ (.A(_2755_),
    .B(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__mux2_1 _6577_ (.A0(_2752_),
    .A1(_2812_),
    .S(_2777_),
    .X(_2813_));
 sky130_fd_sc_hd__inv_2 _6578_ (.A(_2813_),
    .Y(_2814_));
 sky130_fd_sc_hd__nor2_1 _6579_ (.A(net153),
    .B(_2813_),
    .Y(_2815_));
 sky130_fd_sc_hd__nand2_1 _6580_ (.A(net153),
    .B(_2813_),
    .Y(_2816_));
 sky130_fd_sc_hd__and2_1 _6581_ (.A(net122),
    .B(net110),
    .X(_2817_));
 sky130_fd_sc_hd__a211o_1 _6582_ (.A1(_2772_),
    .A2(_2776_),
    .B1(_2817_),
    .C1(_2755_),
    .X(_2818_));
 sky130_fd_sc_hd__nand3b_1 _6583_ (.A_N(net122),
    .B(_2772_),
    .C(_2776_),
    .Y(_2819_));
 sky130_fd_sc_hd__nand2_1 _6584_ (.A(_2818_),
    .B(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__inv_2 _6585_ (.A(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__and3_1 _6586_ (.A(net109),
    .B(_2818_),
    .C(_2819_),
    .X(_2822_));
 sky130_fd_sc_hd__a21oi_2 _6587_ (.A1(_2818_),
    .A2(_2819_),
    .B1(net109),
    .Y(_2823_));
 sky130_fd_sc_hd__nor2_1 _6588_ (.A(net125),
    .B(net110),
    .Y(_2824_));
 sky130_fd_sc_hd__o21bai_4 _6589_ (.A1(_2823_),
    .A2(_2824_),
    .B1_N(_2822_),
    .Y(_2825_));
 sky130_fd_sc_hd__a21oi_4 _6590_ (.A1(_2816_),
    .A2(_2825_),
    .B1(_2815_),
    .Y(_2826_));
 sky130_fd_sc_hd__o21ba_1 _6591_ (.A1(_2810_),
    .A2(_2826_),
    .B1_N(_2808_),
    .X(_2827_));
 sky130_fd_sc_hd__nand2b_1 _6592_ (.A_N(_2804_),
    .B(_2808_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor2_1 _6593_ (.A(_2803_),
    .B(_2804_),
    .Y(_2829_));
 sky130_fd_sc_hd__o311ai_4 _6594_ (.A1(_2804_),
    .A2(_2810_),
    .A3(_2826_),
    .B1(_2828_),
    .C1(_2802_),
    .Y(_2830_));
 sky130_fd_sc_hd__a21o_1 _6595_ (.A1(_2797_),
    .A2(_2830_),
    .B1(_2796_),
    .X(_2831_));
 sky130_fd_sc_hd__and2_1 _6596_ (.A(_2792_),
    .B(_2796_),
    .X(_2832_));
 sky130_fd_sc_hd__and2_1 _6597_ (.A(_2790_),
    .B(_2792_),
    .X(_2833_));
 sky130_fd_sc_hd__a311o_1 _6598_ (.A1(_2792_),
    .A2(_2797_),
    .A3(_2830_),
    .B1(_2832_),
    .C1(_2791_),
    .X(_2834_));
 sky130_fd_sc_hd__nand2_1 _6599_ (.A(net138),
    .B(_2782_),
    .Y(_2835_));
 sky130_fd_sc_hd__and2_1 _6600_ (.A(_2783_),
    .B(_2835_),
    .X(_2836_));
 sky130_fd_sc_hd__nand2_1 _6601_ (.A(net230),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__a211o_4 _6602_ (.A1(_2834_),
    .A2(_2836_),
    .B1(_2780_),
    .C1(_2784_),
    .X(_2838_));
 sky130_fd_sc_hd__xor2_1 _6603_ (.A(_2797_),
    .B(_2830_),
    .X(_2839_));
 sky130_fd_sc_hd__mux2_2 _6604_ (.A0(_2795_),
    .A1(_2839_),
    .S(_2838_),
    .X(_2840_));
 sky130_fd_sc_hd__and2_1 _6605_ (.A(_3477_),
    .B(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__xnor2_2 _6606_ (.A(net140),
    .B(_2840_),
    .Y(_2842_));
 sky130_fd_sc_hd__xor2_1 _6607_ (.A(_2827_),
    .B(_2829_),
    .X(_2843_));
 sky130_fd_sc_hd__xnor2_1 _6608_ (.A(_2827_),
    .B(_2829_),
    .Y(_2844_));
 sky130_fd_sc_hd__mux2_4 _6609_ (.A0(_2801_),
    .A1(_2844_),
    .S(_2838_),
    .X(_2845_));
 sky130_fd_sc_hd__mux2_1 _6610_ (.A0(_2800_),
    .A1(_2843_),
    .S(net227),
    .X(_2846_));
 sky130_fd_sc_hd__nor2_1 _6611_ (.A(net244),
    .B(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nor2_1 _6612_ (.A(_3476_),
    .B(_2845_),
    .Y(_2848_));
 sky130_fd_sc_hd__xnor2_1 _6613_ (.A(_2809_),
    .B(_2826_),
    .Y(_2849_));
 sky130_fd_sc_hd__mux2_2 _6614_ (.A0(_2807_),
    .A1(_2849_),
    .S(_2838_),
    .X(_2850_));
 sky130_fd_sc_hd__and2_1 _6615_ (.A(_3475_),
    .B(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__o211a_1 _6616_ (.A1(_3476_),
    .A2(_2845_),
    .B1(_2850_),
    .C1(_3475_),
    .X(_2852_));
 sky130_fd_sc_hd__nor2_1 _6617_ (.A(_2847_),
    .B(_2848_),
    .Y(_2853_));
 sky130_fd_sc_hd__and2b_1 _6618_ (.A_N(_2815_),
    .B(_2816_),
    .X(_2854_));
 sky130_fd_sc_hd__xor2_1 _6619_ (.A(_2825_),
    .B(_2854_),
    .X(_2855_));
 sky130_fd_sc_hd__mux2_2 _6620_ (.A0(_2814_),
    .A1(_2855_),
    .S(_2838_),
    .X(_2856_));
 sky130_fd_sc_hd__nor2_1 _6621_ (.A(_2822_),
    .B(_2823_),
    .Y(_2857_));
 sky130_fd_sc_hd__xnor2_1 _6622_ (.A(_2824_),
    .B(_2857_),
    .Y(_2858_));
 sky130_fd_sc_hd__mux2_2 _6623_ (.A0(_2821_),
    .A1(_2858_),
    .S(_2838_),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_1 _6624_ (.A(net107),
    .B(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__xnor2_2 _6625_ (.A(net153),
    .B(_2859_),
    .Y(_2861_));
 sky130_fd_sc_hd__nand2_1 _6626_ (.A(net125),
    .B(net110),
    .Y(_2862_));
 sky130_fd_sc_hd__nand3b_1 _6627_ (.A_N(_2824_),
    .B(net227),
    .C(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__or2_1 _6628_ (.A(net125),
    .B(net227),
    .X(_2864_));
 sky130_fd_sc_hd__and3_1 _6629_ (.A(net109),
    .B(_2863_),
    .C(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__nand2_1 _6630_ (.A(_3434_),
    .B(net158),
    .Y(_2866_));
 sky130_fd_sc_hd__a21o_1 _6631_ (.A1(_2863_),
    .A2(_2864_),
    .B1(net109),
    .X(_2867_));
 sky130_fd_sc_hd__and2b_1 _6632_ (.A_N(_2865_),
    .B(_2867_),
    .X(_2868_));
 sky130_fd_sc_hd__a21o_1 _6633_ (.A1(_2866_),
    .A2(_2867_),
    .B1(_2865_),
    .X(_2869_));
 sky130_fd_sc_hd__a21bo_1 _6634_ (.A1(_2861_),
    .A2(_2869_),
    .B1_N(_2860_),
    .X(_2870_));
 sky130_fd_sc_hd__a22o_1 _6635_ (.A1(net106),
    .A2(_2856_),
    .B1(_2859_),
    .B2(net107),
    .X(_2871_));
 sky130_fd_sc_hd__o21a_1 _6636_ (.A1(net106),
    .A2(_2856_),
    .B1(_2871_),
    .X(_2872_));
 sky130_fd_sc_hd__xnor2_1 _6637_ (.A(net150),
    .B(_2856_),
    .Y(_2873_));
 sky130_fd_sc_hd__a31o_4 _6638_ (.A1(_2861_),
    .A2(_2869_),
    .A3(_2873_),
    .B1(_2872_),
    .X(_2874_));
 sky130_fd_sc_hd__nor2_1 _6639_ (.A(_3475_),
    .B(_2850_),
    .Y(_2875_));
 sky130_fd_sc_hd__nor2_2 _6640_ (.A(_2851_),
    .B(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__a311o_1 _6641_ (.A1(_2853_),
    .A2(_2874_),
    .A3(_2876_),
    .B1(_2852_),
    .C1(_2847_),
    .X(_2877_));
 sky130_fd_sc_hd__nor2_1 _6642_ (.A(_2842_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__xnor2_1 _6643_ (.A(_2831_),
    .B(_2833_),
    .Y(_2879_));
 sky130_fd_sc_hd__mux2_2 _6644_ (.A0(_2789_),
    .A1(_2879_),
    .S(_2838_),
    .X(_2880_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(net137),
    .B(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__nor2_1 _6646_ (.A(net137),
    .B(_2880_),
    .Y(_2882_));
 sky130_fd_sc_hd__xnor2_2 _6647_ (.A(_3478_),
    .B(_2880_),
    .Y(_2883_));
 sky130_fd_sc_hd__and4_2 _6648_ (.A(_2842_),
    .B(_2853_),
    .C(_2876_),
    .D(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__o211a_1 _6649_ (.A1(_2847_),
    .A2(_2852_),
    .B1(_2883_),
    .C1(_2842_),
    .X(_2885_));
 sky130_fd_sc_hd__a21o_1 _6650_ (.A1(_2841_),
    .A2(_2881_),
    .B1(_2882_),
    .X(_2886_));
 sky130_fd_sc_hd__or2_1 _6651_ (.A(_2834_),
    .B(_2836_),
    .X(_2887_));
 sky130_fd_sc_hd__nor2_1 _6652_ (.A(_2782_),
    .B(net227),
    .Y(_2888_));
 sky130_fd_sc_hd__a31oi_1 _6653_ (.A1(_2837_),
    .A2(net227),
    .A3(_2887_),
    .B1(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__a21oi_1 _6654_ (.A1(_2783_),
    .A2(_2837_),
    .B1(_2779_),
    .Y(_2890_));
 sky130_fd_sc_hd__a21o_1 _6655_ (.A1(_2772_),
    .A2(_2773_),
    .B1(_2775_),
    .X(_2891_));
 sky130_fd_sc_hd__nand2_1 _6656_ (.A(_1797_),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__or3b_4 _6657_ (.A(_2892_),
    .B(_2890_),
    .C_N(_2889_),
    .X(_2893_));
 sky130_fd_sc_hd__or3_4 _6658_ (.A(_2885_),
    .B(_2886_),
    .C(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__a21oi_4 _6659_ (.A1(net236),
    .A2(_2884_),
    .B1(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__a21o_4 _6660_ (.A1(_2874_),
    .A2(_2884_),
    .B1(_2894_),
    .X(_2896_));
 sky130_fd_sc_hd__a21o_1 _6661_ (.A1(_2842_),
    .A2(_2877_),
    .B1(_2895_),
    .X(_2897_));
 sky130_fd_sc_hd__o2bb2a_4 _6662_ (.A1_N(_2840_),
    .A2_N(_2895_),
    .B1(_2897_),
    .B2(_2878_),
    .X(_2898_));
 sky130_fd_sc_hd__and2_4 _6663_ (.A(net137),
    .B(_2898_),
    .X(_2899_));
 sky130_fd_sc_hd__nand2_1 _6664_ (.A(net137),
    .B(_2898_),
    .Y(_2900_));
 sky130_fd_sc_hd__a21o_1 _6665_ (.A1(_2874_),
    .A2(_2876_),
    .B1(_2851_),
    .X(_2901_));
 sky130_fd_sc_hd__xnor2_1 _6666_ (.A(_2853_),
    .B(_2901_),
    .Y(_2902_));
 sky130_fd_sc_hd__mux2_2 _6667_ (.A0(_2846_),
    .A1(_2902_),
    .S(_2896_),
    .X(_2903_));
 sky130_fd_sc_hd__and2_1 _6668_ (.A(net140),
    .B(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__xnor2_1 _6669_ (.A(net140),
    .B(_2903_),
    .Y(_2905_));
 sky130_fd_sc_hd__xor2_1 _6670_ (.A(_2874_),
    .B(_2876_),
    .X(_2906_));
 sky130_fd_sc_hd__mux2_2 _6671_ (.A0(_2850_),
    .A1(_2906_),
    .S(_2896_),
    .X(_2907_));
 sky130_fd_sc_hd__and2_1 _6672_ (.A(_3476_),
    .B(_2907_),
    .X(_2908_));
 sky130_fd_sc_hd__nor2_1 _6673_ (.A(_3476_),
    .B(_2907_),
    .Y(_2909_));
 sky130_fd_sc_hd__nor2_2 _6674_ (.A(_2908_),
    .B(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__and2b_1 _6675_ (.A_N(_2905_),
    .B(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__xnor2_1 _6676_ (.A(_2866_),
    .B(_2868_),
    .Y(_2912_));
 sky130_fd_sc_hd__a221o_1 _6677_ (.A1(_2863_),
    .A2(_2864_),
    .B1(_2874_),
    .B2(_2884_),
    .C1(_2894_),
    .X(_2913_));
 sky130_fd_sc_hd__a21bo_1 _6678_ (.A1(_2896_),
    .A2(_2912_),
    .B1_N(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__inv_2 _6679_ (.A(_2914_),
    .Y(_2915_));
 sky130_fd_sc_hd__nor2_1 _6680_ (.A(net153),
    .B(_2914_),
    .Y(_2916_));
 sky130_fd_sc_hd__nand2_1 _6681_ (.A(net153),
    .B(_2914_),
    .Y(_2917_));
 sky130_fd_sc_hd__a211o_1 _6682_ (.A1(net236),
    .A2(_2884_),
    .B1(_2894_),
    .C1(net128),
    .X(_2918_));
 sky130_fd_sc_hd__nand2_1 _6683_ (.A(net128),
    .B(net110),
    .Y(_2919_));
 sky130_fd_sc_hd__and2_1 _6684_ (.A(_2866_),
    .B(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__nand2_1 _6685_ (.A(_2866_),
    .B(_2919_),
    .Y(_2921_));
 sky130_fd_sc_hd__a211o_1 _6686_ (.A1(net236),
    .A2(_2884_),
    .B1(_2894_),
    .C1(_3434_),
    .X(_2922_));
 sky130_fd_sc_hd__o21a_1 _6687_ (.A1(_2895_),
    .A2(_2921_),
    .B1(_2918_),
    .X(_2923_));
 sky130_fd_sc_hd__o211a_1 _6688_ (.A1(_2895_),
    .A2(_2921_),
    .B1(_2918_),
    .C1(net109),
    .X(_2924_));
 sky130_fd_sc_hd__o211ai_1 _6689_ (.A1(_2895_),
    .A2(_2920_),
    .B1(_2922_),
    .C1(net156),
    .Y(_2925_));
 sky130_fd_sc_hd__xor2_1 _6690_ (.A(net129),
    .B(net158),
    .X(_2926_));
 sky130_fd_sc_hd__nand2_1 _6691_ (.A(_3435_),
    .B(net158),
    .Y(_2927_));
 sky130_fd_sc_hd__a21o_1 _6692_ (.A1(_2925_),
    .A2(_2927_),
    .B1(_2924_),
    .X(_2928_));
 sky130_fd_sc_hd__a21o_1 _6693_ (.A1(_2917_),
    .A2(_2928_),
    .B1(_2916_),
    .X(_2929_));
 sky130_fd_sc_hd__xor2_1 _6694_ (.A(_2861_),
    .B(_2869_),
    .X(_2930_));
 sky130_fd_sc_hd__mux2_4 _6695_ (.A0(_2859_),
    .A1(_2930_),
    .S(_2896_),
    .X(_2931_));
 sky130_fd_sc_hd__and2_1 _6696_ (.A(net106),
    .B(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__nor2_1 _6697_ (.A(net106),
    .B(_2931_),
    .Y(_2933_));
 sky130_fd_sc_hd__nor2_2 _6698_ (.A(_2932_),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__xor2_1 _6699_ (.A(_2870_),
    .B(_2873_),
    .X(_2935_));
 sky130_fd_sc_hd__mux2_4 _6700_ (.A0(_2856_),
    .A1(_2935_),
    .S(_2896_),
    .X(_2936_));
 sky130_fd_sc_hd__inv_2 _6701_ (.A(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hd__xnor2_1 _6702_ (.A(net147),
    .B(_2936_),
    .Y(_2938_));
 sky130_fd_sc_hd__o211a_1 _6703_ (.A1(_3475_),
    .A2(_2936_),
    .B1(_2931_),
    .C1(net106),
    .X(_2939_));
 sky130_fd_sc_hd__a21o_1 _6704_ (.A1(_3475_),
    .A2(_2936_),
    .B1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__a31o_4 _6705_ (.A1(_2929_),
    .A2(_2934_),
    .A3(_2938_),
    .B1(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__o21ba_4 _6706_ (.A1(net140),
    .A2(_2903_),
    .B1_N(_2908_),
    .X(_2942_));
 sky130_fd_sc_hd__a21o_1 _6707_ (.A1(_2842_),
    .A2(_2877_),
    .B1(_2841_),
    .X(_2943_));
 sky130_fd_sc_hd__xnor2_1 _6708_ (.A(_2883_),
    .B(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__mux2_1 _6709_ (.A0(_2880_),
    .A1(_2944_),
    .S(_2896_),
    .X(_2945_));
 sky130_fd_sc_hd__or2_4 _6710_ (.A(net138),
    .B(_2898_),
    .X(_2946_));
 sky130_fd_sc_hd__o311ai_4 _6711_ (.A1(_2899_),
    .A2(_2904_),
    .A3(_2942_),
    .B1(_2945_),
    .C1(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__a31o_4 _6712_ (.A1(_2900_),
    .A2(_2911_),
    .A3(_2941_),
    .B1(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__a21o_1 _6713_ (.A1(_2929_),
    .A2(_2934_),
    .B1(_2932_),
    .X(_2949_));
 sky130_fd_sc_hd__xnor2_1 _6714_ (.A(_2938_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__mux2_2 _6715_ (.A0(_2937_),
    .A1(_2950_),
    .S(_2948_),
    .X(_2951_));
 sky130_fd_sc_hd__nor2_1 _6716_ (.A(net245),
    .B(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__nand2_1 _6717_ (.A(net144),
    .B(_2951_),
    .Y(_2953_));
 sky130_fd_sc_hd__xnor2_2 _6718_ (.A(net144),
    .B(_2951_),
    .Y(_2954_));
 sky130_fd_sc_hd__xor2_1 _6719_ (.A(_2929_),
    .B(_2934_),
    .X(_2955_));
 sky130_fd_sc_hd__mux2_2 _6720_ (.A0(_2931_),
    .A1(_2955_),
    .S(_2948_),
    .X(_2956_));
 sky130_fd_sc_hd__nand2_1 _6721_ (.A(_3475_),
    .B(_2956_),
    .Y(_2957_));
 sky130_fd_sc_hd__xnor2_4 _6722_ (.A(_3475_),
    .B(_2956_),
    .Y(_2958_));
 sky130_fd_sc_hd__nand2b_1 _6723_ (.A_N(_2916_),
    .B(_2917_),
    .Y(_2959_));
 sky130_fd_sc_hd__xnor2_1 _6724_ (.A(_2928_),
    .B(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__mux2_2 _6725_ (.A0(_2915_),
    .A1(_2960_),
    .S(_2948_),
    .X(_2961_));
 sky130_fd_sc_hd__inv_2 _6726_ (.A(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__nand2_1 _6727_ (.A(net106),
    .B(_2961_),
    .Y(_2963_));
 sky130_fd_sc_hd__nand2b_1 _6728_ (.A_N(_2924_),
    .B(_2925_),
    .Y(_2964_));
 sky130_fd_sc_hd__xnor2_1 _6729_ (.A(_2927_),
    .B(_2964_),
    .Y(_2965_));
 sky130_fd_sc_hd__mux2_4 _6730_ (.A0(_2923_),
    .A1(_2965_),
    .S(_2948_),
    .X(_2966_));
 sky130_fd_sc_hd__inv_2 _6731_ (.A(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__nor2_1 _6732_ (.A(net153),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__o211ai_1 _6733_ (.A1(net106),
    .A2(_2961_),
    .B1(_2966_),
    .C1(net107),
    .Y(_2969_));
 sky130_fd_sc_hd__and2_1 _6734_ (.A(_2963_),
    .B(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__xnor2_2 _6735_ (.A(net106),
    .B(_2961_),
    .Y(_2971_));
 sky130_fd_sc_hd__mux2_4 _6736_ (.A0(net129),
    .A1(_2926_),
    .S(_2948_),
    .X(_2972_));
 sky130_fd_sc_hd__and2_1 _6737_ (.A(net108),
    .B(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__nand2_1 _6738_ (.A(_3436_),
    .B(net158),
    .Y(_2974_));
 sky130_fd_sc_hd__or2_4 _6739_ (.A(net108),
    .B(_2972_),
    .X(_2975_));
 sky130_fd_sc_hd__and2b_1 _6740_ (.A_N(_2973_),
    .B(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__a21o_4 _6741_ (.A1(_2974_),
    .A2(_2975_),
    .B1(_2973_),
    .X(_2977_));
 sky130_fd_sc_hd__xnor2_2 _6742_ (.A(net153),
    .B(_2966_),
    .Y(_2978_));
 sky130_fd_sc_hd__nand3b_1 _6743_ (.A_N(_2971_),
    .B(_2977_),
    .C(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__a21o_1 _6744_ (.A1(_2970_),
    .A2(_2979_),
    .B1(_2958_),
    .X(_2980_));
 sky130_fd_sc_hd__a21oi_1 _6745_ (.A1(_2957_),
    .A2(_2980_),
    .B1(_2954_),
    .Y(_2981_));
 sky130_fd_sc_hd__a21oi_1 _6746_ (.A1(_2910_),
    .A2(_2941_),
    .B1(_2908_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _6747_ (.A(_2905_),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__o21a_1 _6748_ (.A1(_2905_),
    .A2(_2982_),
    .B1(net225),
    .X(_2984_));
 sky130_fd_sc_hd__o2bb2a_2 _6749_ (.A1_N(_2984_),
    .A2_N(_2983_),
    .B1(net225),
    .B2(_2903_),
    .X(_2985_));
 sky130_fd_sc_hd__nand2_1 _6750_ (.A(net137),
    .B(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__xnor2_1 _6751_ (.A(_2910_),
    .B(_2941_),
    .Y(_2987_));
 sky130_fd_sc_hd__a311o_1 _6752_ (.A1(_2900_),
    .A2(_2911_),
    .A3(_2941_),
    .B1(_2947_),
    .C1(_2907_),
    .X(_2988_));
 sky130_fd_sc_hd__a21boi_2 _6753_ (.A1(net225),
    .A2(_2987_),
    .B1_N(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__nand2_1 _6754_ (.A(_3477_),
    .B(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__o21ai_1 _6755_ (.A1(net137),
    .A2(_2985_),
    .B1(_2990_),
    .Y(_2991_));
 sky130_fd_sc_hd__nand2_1 _6756_ (.A(_2900_),
    .B(_2946_),
    .Y(_2992_));
 sky130_fd_sc_hd__o2bb2a_1 _6757_ (.A1_N(_2911_),
    .A2_N(_2941_),
    .B1(_2942_),
    .B2(_2904_),
    .X(_2993_));
 sky130_fd_sc_hd__o21a_1 _6758_ (.A1(_2992_),
    .A2(_2993_),
    .B1(_2948_),
    .X(_2994_));
 sky130_fd_sc_hd__nand2_1 _6759_ (.A(_2992_),
    .B(_2993_),
    .Y(_2995_));
 sky130_fd_sc_hd__a2bb2o_1 _6760_ (.A1_N(_2898_),
    .A2_N(net225),
    .B1(_2994_),
    .B2(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__a21oi_1 _6761_ (.A1(_2946_),
    .A2(_2994_),
    .B1(_2945_),
    .Y(_2997_));
 sky130_fd_sc_hd__a211o_1 _6762_ (.A1(net236),
    .A2(_2884_),
    .B1(_2885_),
    .C1(_2886_),
    .X(_2998_));
 sky130_fd_sc_hd__nand2b_1 _6763_ (.A_N(_2889_),
    .B(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__or4b_4 _6764_ (.A(_2890_),
    .B(_2892_),
    .C(_2997_),
    .D_N(_2999_),
    .X(_3000_));
 sky130_fd_sc_hd__a211o_4 _6765_ (.A1(_2986_),
    .A2(_2991_),
    .B1(_2996_),
    .C1(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__nor4b_4 _6766_ (.A(_2954_),
    .B(_2958_),
    .C(_2971_),
    .D_N(_2978_),
    .Y(_3002_));
 sky130_fd_sc_hd__a211oi_1 _6767_ (.A1(_2963_),
    .A2(_2969_),
    .B1(_2954_),
    .C1(_2958_),
    .Y(_3003_));
 sky130_fd_sc_hd__a31o_1 _6768_ (.A1(_3475_),
    .A2(_2953_),
    .A3(_2956_),
    .B1(_2952_),
    .X(_3004_));
 sky130_fd_sc_hd__a211oi_1 _6769_ (.A1(_2977_),
    .A2(_3002_),
    .B1(_3003_),
    .C1(_3004_),
    .Y(_3005_));
 sky130_fd_sc_hd__a211o_4 _6770_ (.A1(_2977_),
    .A2(_3002_),
    .B1(_3003_),
    .C1(_3004_),
    .X(_3006_));
 sky130_fd_sc_hd__xnor2_1 _6771_ (.A(net140),
    .B(_2989_),
    .Y(_3007_));
 sky130_fd_sc_hd__inv_2 _6772_ (.A(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__xnor2_2 _6773_ (.A(net137),
    .B(_2985_),
    .Y(_3009_));
 sky130_fd_sc_hd__nor2_2 _6774_ (.A(_3008_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__a21oi_2 _6775_ (.A1(_3006_),
    .A2(_3010_),
    .B1(_3001_),
    .Y(_3011_));
 sky130_fd_sc_hd__a21o_4 _6776_ (.A1(_3006_),
    .A2(_3010_),
    .B1(_3001_),
    .X(_3012_));
 sky130_fd_sc_hd__a31o_1 _6777_ (.A1(_2954_),
    .A2(_2957_),
    .A3(_2980_),
    .B1(_3011_),
    .X(_3013_));
 sky130_fd_sc_hd__o22a_2 _6778_ (.A1(_2951_),
    .A2(net243),
    .B1(_3013_),
    .B2(_2981_),
    .X(_3014_));
 sky130_fd_sc_hd__inv_2 _6779_ (.A(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__or2_1 _6780_ (.A(net142),
    .B(_3014_),
    .X(_3016_));
 sky130_fd_sc_hd__nand3_1 _6781_ (.A(_2958_),
    .B(_2970_),
    .C(_2979_),
    .Y(_3017_));
 sky130_fd_sc_hd__and3_1 _6782_ (.A(_2980_),
    .B(_3012_),
    .C(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__a21oi_2 _6783_ (.A1(_2956_),
    .A2(_3011_),
    .B1(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__xnor2_1 _6784_ (.A(net145),
    .B(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__a21oi_1 _6785_ (.A1(_2977_),
    .A2(_2978_),
    .B1(_2968_),
    .Y(_3021_));
 sky130_fd_sc_hd__xnor2_1 _6786_ (.A(_2971_),
    .B(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__mux2_1 _6787_ (.A0(_2962_),
    .A1(_3022_),
    .S(_3012_),
    .X(_3023_));
 sky130_fd_sc_hd__and2_1 _6788_ (.A(net148),
    .B(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__xnor2_1 _6789_ (.A(_2977_),
    .B(_2978_),
    .Y(_3025_));
 sky130_fd_sc_hd__mux2_4 _6790_ (.A0(_2967_),
    .A1(_3025_),
    .S(_3012_),
    .X(_3026_));
 sky130_fd_sc_hd__inv_2 _6791_ (.A(_3026_),
    .Y(_3027_));
 sky130_fd_sc_hd__nor2_1 _6792_ (.A(net151),
    .B(_3026_),
    .Y(_3028_));
 sky130_fd_sc_hd__nor2_1 _6793_ (.A(net148),
    .B(_3023_),
    .Y(_3029_));
 sky130_fd_sc_hd__o22a_1 _6794_ (.A1(net147),
    .A2(_3023_),
    .B1(_3026_),
    .B2(net151),
    .X(_3030_));
 sky130_fd_sc_hd__xnor2_4 _6795_ (.A(net151),
    .B(_3026_),
    .Y(_3031_));
 sky130_fd_sc_hd__xnor2_1 _6796_ (.A(_2974_),
    .B(_2976_),
    .Y(_3032_));
 sky130_fd_sc_hd__a211oi_1 _6797_ (.A1(net231),
    .A2(_3010_),
    .B1(_2972_),
    .C1(_3001_),
    .Y(_3033_));
 sky130_fd_sc_hd__a21o_1 _6798_ (.A1(_3012_),
    .A2(_3032_),
    .B1(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__and2_1 _6799_ (.A(net154),
    .B(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__a211o_1 _6800_ (.A1(_3012_),
    .A2(_3032_),
    .B1(_3033_),
    .C1(net154),
    .X(_3036_));
 sky130_fd_sc_hd__a211oi_2 _6801_ (.A1(net232),
    .A2(_3010_),
    .B1(net131),
    .C1(_3001_),
    .Y(_3037_));
 sky130_fd_sc_hd__xnor2_2 _6802_ (.A(net131),
    .B(net158),
    .Y(_3038_));
 sky130_fd_sc_hd__a211o_1 _6803_ (.A1(net231),
    .A2(_3010_),
    .B1(_3436_),
    .C1(_3001_),
    .X(_3039_));
 sky130_fd_sc_hd__a21oi_2 _6804_ (.A1(net243),
    .A2(_3038_),
    .B1(_3037_),
    .Y(_3040_));
 sky130_fd_sc_hd__a211o_1 _6805_ (.A1(_3012_),
    .A2(_3038_),
    .B1(_3037_),
    .C1(net156),
    .X(_3041_));
 sky130_fd_sc_hd__o211a_1 _6806_ (.A1(_3011_),
    .A2(_3038_),
    .B1(_3039_),
    .C1(net156),
    .X(_3042_));
 sky130_fd_sc_hd__xnor2_1 _6807_ (.A(net157),
    .B(_3040_),
    .Y(_3043_));
 sky130_fd_sc_hd__nor2_1 _6808_ (.A(net134),
    .B(net111),
    .Y(_3044_));
 sky130_fd_sc_hd__inv_2 _6809_ (.A(_3044_),
    .Y(_3045_));
 sky130_fd_sc_hd__nand2_1 _6810_ (.A(_3043_),
    .B(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__and2_1 _6811_ (.A(_3041_),
    .B(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__o211a_1 _6812_ (.A1(_3042_),
    .A2(_3044_),
    .B1(_3036_),
    .C1(_3041_),
    .X(_3048_));
 sky130_fd_sc_hd__nor3_1 _6813_ (.A(_3031_),
    .B(_3035_),
    .C(_3048_),
    .Y(_3049_));
 sky130_fd_sc_hd__o31a_1 _6814_ (.A1(_3031_),
    .A2(_3035_),
    .A3(_3048_),
    .B1(_3030_),
    .X(_3050_));
 sky130_fd_sc_hd__or2_1 _6815_ (.A(_3024_),
    .B(_3029_),
    .X(_3051_));
 sky130_fd_sc_hd__nor2_1 _6816_ (.A(_3024_),
    .B(_3050_),
    .Y(_3052_));
 sky130_fd_sc_hd__or3_1 _6817_ (.A(_3020_),
    .B(_3024_),
    .C(_3050_),
    .X(_3053_));
 sky130_fd_sc_hd__o21ai_1 _6818_ (.A1(net145),
    .A2(_3019_),
    .B1(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__a211o_1 _6819_ (.A1(net142),
    .A2(_3014_),
    .B1(_3019_),
    .C1(net242),
    .X(_3055_));
 sky130_fd_sc_hd__xnor2_1 _6820_ (.A(net142),
    .B(_3014_),
    .Y(_3056_));
 sky130_fd_sc_hd__o41a_1 _6821_ (.A1(_3020_),
    .A2(_3024_),
    .A3(_3050_),
    .A4(_3056_),
    .B1(_3055_),
    .X(_3057_));
 sky130_fd_sc_hd__nand2_1 _6822_ (.A(_3006_),
    .B(_3007_),
    .Y(_3058_));
 sky130_fd_sc_hd__nand2_1 _6823_ (.A(_3005_),
    .B(_3008_),
    .Y(_3059_));
 sky130_fd_sc_hd__and3_1 _6824_ (.A(net243),
    .B(_3058_),
    .C(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__a21oi_1 _6825_ (.A1(_2989_),
    .A2(_3011_),
    .B1(_3060_),
    .Y(_3061_));
 sky130_fd_sc_hd__or2_1 _6826_ (.A(net139),
    .B(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__nand2_1 _6827_ (.A(net139),
    .B(_3061_),
    .Y(_3063_));
 sky130_fd_sc_hd__nand2_1 _6828_ (.A(_3062_),
    .B(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__a21o_2 _6829_ (.A1(_3016_),
    .A2(_3057_),
    .B1(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__a21o_1 _6830_ (.A1(_2990_),
    .A2(_3058_),
    .B1(_3009_),
    .X(_3066_));
 sky130_fd_sc_hd__and3_1 _6831_ (.A(_2990_),
    .B(_3009_),
    .C(_3058_),
    .X(_3067_));
 sky130_fd_sc_hd__nand2_1 _6832_ (.A(net243),
    .B(_3066_),
    .Y(_3068_));
 sky130_fd_sc_hd__o22a_1 _6833_ (.A1(_2985_),
    .A2(net243),
    .B1(_3067_),
    .B2(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__a22o_1 _6834_ (.A1(_2986_),
    .A2(_2991_),
    .B1(_3006_),
    .B2(_3010_),
    .X(_3070_));
 sky130_fd_sc_hd__a21o_1 _6835_ (.A1(_2996_),
    .A2(_3070_),
    .B1(_3000_),
    .X(_3071_));
 sky130_fd_sc_hd__and3b_2 _6836_ (.A_N(_3071_),
    .B(_3062_),
    .C(_3069_),
    .X(_3072_));
 sky130_fd_sc_hd__nand2_4 _6837_ (.A(_3065_),
    .B(_3072_),
    .Y(_3073_));
 sky130_fd_sc_hd__xnor2_1 _6838_ (.A(_3054_),
    .B(_3056_),
    .Y(_3074_));
 sky130_fd_sc_hd__mux2_2 _6839_ (.A0(_3015_),
    .A1(_3074_),
    .S(_3073_),
    .X(_3075_));
 sky130_fd_sc_hd__xnor2_2 _6840_ (.A(_3478_),
    .B(_3075_),
    .Y(_3076_));
 sky130_fd_sc_hd__xor2_1 _6841_ (.A(_3020_),
    .B(_3052_),
    .X(_3077_));
 sky130_fd_sc_hd__mux2_1 _6842_ (.A0(_3019_),
    .A1(_3077_),
    .S(_3073_),
    .X(_3078_));
 sky130_fd_sc_hd__nor2_1 _6843_ (.A(net142),
    .B(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__and2_1 _6844_ (.A(net142),
    .B(_3078_),
    .X(_3080_));
 sky130_fd_sc_hd__nor2_1 _6845_ (.A(_3079_),
    .B(_3080_),
    .Y(_3081_));
 sky130_fd_sc_hd__inv_2 _6846_ (.A(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__o21ai_1 _6847_ (.A1(_3028_),
    .A2(_3049_),
    .B1(_3051_),
    .Y(_3083_));
 sky130_fd_sc_hd__or3_1 _6848_ (.A(_3028_),
    .B(_3049_),
    .C(_3051_),
    .X(_3084_));
 sky130_fd_sc_hd__a22o_1 _6849_ (.A1(_3065_),
    .A2(_3072_),
    .B1(_3083_),
    .B2(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__o21a_1 _6850_ (.A1(_3023_),
    .A2(_3073_),
    .B1(_3085_),
    .X(_3086_));
 sky130_fd_sc_hd__and2_1 _6851_ (.A(net145),
    .B(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__nand2_1 _6852_ (.A(net238),
    .B(_3086_),
    .Y(_3088_));
 sky130_fd_sc_hd__o21a_1 _6853_ (.A1(_3035_),
    .A2(_3048_),
    .B1(_3031_),
    .X(_3089_));
 sky130_fd_sc_hd__nor2_1 _6854_ (.A(_3049_),
    .B(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__mux2_1 _6855_ (.A0(_3027_),
    .A1(_3090_),
    .S(_3073_),
    .X(_3091_));
 sky130_fd_sc_hd__and2_1 _6856_ (.A(_3475_),
    .B(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__xnor2_1 _6857_ (.A(_3475_),
    .B(_3091_),
    .Y(_3093_));
 sky130_fd_sc_hd__inv_2 _6858_ (.A(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__and2b_1 _6859_ (.A_N(_3035_),
    .B(_3036_),
    .X(_3095_));
 sky130_fd_sc_hd__xor2_1 _6860_ (.A(_3047_),
    .B(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__a21o_1 _6861_ (.A1(_3065_),
    .A2(_3072_),
    .B1(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__nand3b_1 _6862_ (.A_N(_3034_),
    .B(_3065_),
    .C(_3072_),
    .Y(_3098_));
 sky130_fd_sc_hd__nand2_1 _6863_ (.A(_3097_),
    .B(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__and3_1 _6864_ (.A(net151),
    .B(_3097_),
    .C(_3098_),
    .X(_3100_));
 sky130_fd_sc_hd__or2_1 _6865_ (.A(_3043_),
    .B(_3045_),
    .X(_3101_));
 sky130_fd_sc_hd__a22o_1 _6866_ (.A1(_3065_),
    .A2(_3072_),
    .B1(_3101_),
    .B2(_3046_),
    .X(_3102_));
 sky130_fd_sc_hd__o21a_1 _6867_ (.A1(_3040_),
    .A2(_3073_),
    .B1(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__o211ai_2 _6868_ (.A1(_3040_),
    .A2(_3073_),
    .B1(_3102_),
    .C1(net107),
    .Y(_3104_));
 sky130_fd_sc_hd__and2_1 _6869_ (.A(net106),
    .B(_3099_),
    .X(_3105_));
 sky130_fd_sc_hd__a21o_1 _6870_ (.A1(_3097_),
    .A2(_3098_),
    .B1(net151),
    .X(_3106_));
 sky130_fd_sc_hd__xnor2_2 _6871_ (.A(net107),
    .B(_3103_),
    .Y(_3107_));
 sky130_fd_sc_hd__or2_1 _6872_ (.A(net133),
    .B(net160),
    .X(_3108_));
 sky130_fd_sc_hd__a22o_1 _6873_ (.A1(net235),
    .A2(_3072_),
    .B1(_3108_),
    .B2(_2098_),
    .X(_3109_));
 sky130_fd_sc_hd__nand3_1 _6874_ (.A(_3437_),
    .B(net235),
    .C(_3072_),
    .Y(_3110_));
 sky130_fd_sc_hd__and3_1 _6875_ (.A(net108),
    .B(_3109_),
    .C(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__a21o_1 _6876_ (.A1(_3109_),
    .A2(_3110_),
    .B1(net108),
    .X(_3112_));
 sky130_fd_sc_hd__and2b_1 _6877_ (.A_N(_3111_),
    .B(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__a21oi_2 _6878_ (.A1(_2519_),
    .A2(_3112_),
    .B1(_3111_),
    .Y(_3114_));
 sky130_fd_sc_hd__a21o_1 _6879_ (.A1(_3104_),
    .A2(_3106_),
    .B1(_3100_),
    .X(_3115_));
 sky130_fd_sc_hd__nor2_1 _6880_ (.A(_3100_),
    .B(_3105_),
    .Y(_3116_));
 sky130_fd_sc_hd__o41ai_4 _6881_ (.A1(_3100_),
    .A2(_3105_),
    .A3(_3107_),
    .A4(_3114_),
    .B1(_3115_),
    .Y(_3117_));
 sky130_fd_sc_hd__nor2_1 _6882_ (.A(net238),
    .B(_3086_),
    .Y(_3118_));
 sky130_fd_sc_hd__a21o_1 _6883_ (.A1(_3088_),
    .A2(_3092_),
    .B1(_3118_),
    .X(_3119_));
 sky130_fd_sc_hd__nor2_1 _6884_ (.A(_3087_),
    .B(_3118_),
    .Y(_3120_));
 sky130_fd_sc_hd__a31o_1 _6885_ (.A1(_3094_),
    .A2(_3117_),
    .A3(_3120_),
    .B1(_3119_),
    .X(_3121_));
 sky130_fd_sc_hd__a31oi_2 _6886_ (.A1(_3094_),
    .A2(_3117_),
    .A3(_3120_),
    .B1(_3119_),
    .Y(_3122_));
 sky130_fd_sc_hd__nand2_1 _6887_ (.A(_3081_),
    .B(_3121_),
    .Y(_3123_));
 sky130_fd_sc_hd__nand2_1 _6888_ (.A(net235),
    .B(_3073_),
    .Y(_3124_));
 sky130_fd_sc_hd__a21oi_1 _6889_ (.A1(_3062_),
    .A2(net235),
    .B1(_3069_),
    .Y(_3125_));
 sky130_fd_sc_hd__a31oi_1 _6890_ (.A1(_3016_),
    .A2(_3057_),
    .A3(_3064_),
    .B1(_3124_),
    .Y(_3126_));
 sky130_fd_sc_hd__nor2_1 _6891_ (.A(_3061_),
    .B(_3073_),
    .Y(_3127_));
 sky130_fd_sc_hd__a2111o_1 _6892_ (.A1(_3478_),
    .A2(_3075_),
    .B1(_3126_),
    .C1(_3127_),
    .D1(_3071_),
    .X(_3128_));
 sky130_fd_sc_hd__nor2_1 _6893_ (.A(_3125_),
    .B(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__o21ai_1 _6894_ (.A1(_3478_),
    .A2(_3075_),
    .B1(_3079_),
    .Y(_3130_));
 sky130_fd_sc_hd__o311a_4 _6895_ (.A1(_3076_),
    .A2(_3082_),
    .A3(_3122_),
    .B1(_3129_),
    .C1(_3130_),
    .X(_3131_));
 sky130_fd_sc_hd__nand2_4 _6896_ (.A(_3131_),
    .B(net162),
    .Y(_3132_));
 sky130_fd_sc_hd__mux2_4 _6897_ (.A0(net135),
    .A1(_2544_),
    .S(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__o211a_1 _6898_ (.A1(net161),
    .A2(_2544_),
    .B1(_3132_),
    .C1(net97),
    .X(_3134_));
 sky130_fd_sc_hd__a21oi_1 _6899_ (.A1(_3505_),
    .A2(_3514_),
    .B1(_2543_),
    .Y(_3135_));
 sky130_fd_sc_hd__nand2_1 _6900_ (.A(net162),
    .B(net101),
    .Y(_3136_));
 sky130_fd_sc_hd__a21oi_1 _6901_ (.A1(_0500_),
    .A2(_3136_),
    .B1(_2558_),
    .Y(_3137_));
 sky130_fd_sc_hd__a311o_1 _6902_ (.A1(net133),
    .A2(net117),
    .A3(_3517_),
    .B1(_0585_),
    .C1(_3135_),
    .X(_3138_));
 sky130_fd_sc_hd__a2111o_1 _6903_ (.A1(_0502_),
    .A2(_3133_),
    .B1(_3134_),
    .C1(_3137_),
    .D1(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__o31a_1 _6904_ (.A1(net135),
    .A2(net160),
    .A3(_0586_),
    .B1(_0579_),
    .X(_3140_));
 sky130_fd_sc_hd__nand2_1 _6905_ (.A(_3139_),
    .B(_3140_),
    .Y(_3141_));
 sky130_fd_sc_hd__a221o_1 _6906_ (.A1(_0420_),
    .A2(_0574_),
    .B1(_2665_),
    .B2(_3141_),
    .C1(net100),
    .X(_3142_));
 sky130_fd_sc_hd__a32o_1 _6907_ (.A1(net871),
    .A2(_3515_),
    .A3(_3563_),
    .B1(_3570_),
    .B2(net127),
    .X(_3143_));
 sky130_fd_sc_hd__a31o_1 _6908_ (.A1(net133),
    .A2(net117),
    .A3(_3517_),
    .B1(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__or2_1 _6909_ (.A(net63),
    .B(_2544_),
    .X(_3145_));
 sky130_fd_sc_hd__and3_1 _6910_ (.A(_3504_),
    .B(_2559_),
    .C(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__nor2_1 _6911_ (.A(net117),
    .B(_3512_),
    .Y(_3147_));
 sky130_fd_sc_hd__o2bb2a_2 _6912_ (.A1_N(_3508_),
    .A2_N(_3563_),
    .B1(_2571_),
    .B2(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__inv_2 _6913_ (.A(_3148_),
    .Y(_3149_));
 sky130_fd_sc_hd__a21oi_1 _6914_ (.A1(_2559_),
    .A2(_3145_),
    .B1(_3513_),
    .Y(_3150_));
 sky130_fd_sc_hd__a21oi_1 _6915_ (.A1(_3148_),
    .A2(_3150_),
    .B1(_3146_),
    .Y(_3151_));
 sky130_fd_sc_hd__o21ai_1 _6916_ (.A1(_3144_),
    .A2(_3151_),
    .B1(net100),
    .Y(_3152_));
 sky130_fd_sc_hd__a21oi_1 _6917_ (.A1(_3142_),
    .A2(_3152_),
    .B1(net103),
    .Y(_3153_));
 sky130_fd_sc_hd__o31a_1 _6918_ (.A1(net161),
    .A2(_3571_),
    .A3(net94),
    .B1(_3524_),
    .X(_3154_));
 sky130_fd_sc_hd__nand2_1 _6919_ (.A(\as1802.instr_latch[7] ),
    .B(_2586_),
    .Y(_3155_));
 sky130_fd_sc_hd__or4_1 _6920_ (.A(net171),
    .B(\as1802.mem_write ),
    .C(\as1802.lda ),
    .D(_3544_),
    .X(_3156_));
 sky130_fd_sc_hd__a2bb2o_1 _6921_ (.A1_N(_3553_),
    .A2_N(_3154_),
    .B1(_0559_),
    .B2(_0511_),
    .X(_3157_));
 sky130_fd_sc_hd__or4_1 _6922_ (.A(net173),
    .B(_3570_),
    .C(net94),
    .D(_0539_),
    .X(_3158_));
 sky130_fd_sc_hd__o32a_1 _6923_ (.A1(net102),
    .A2(_0534_),
    .A3(_0581_),
    .B1(_3158_),
    .B2(net167),
    .X(_3159_));
 sky130_fd_sc_hd__o2111a_1 _6924_ (.A1(_3553_),
    .A2(_3155_),
    .B1(_3156_),
    .C1(_3557_),
    .D1(_0562_),
    .X(_3160_));
 sky130_fd_sc_hd__and4_1 _6925_ (.A(_2287_),
    .B(_2293_),
    .C(_3159_),
    .D(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__nor3b_4 _6926_ (.A(_2623_),
    .B(_3157_),
    .C_N(_3161_),
    .Y(_3162_));
 sky130_fd_sc_hd__or3b_4 _6927_ (.A(_2623_),
    .B(_3157_),
    .C_N(_3161_),
    .X(_3163_));
 sky130_fd_sc_hd__a21o_1 _6928_ (.A1(net31),
    .A2(net103),
    .B1(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__o221a_1 _6929_ (.A1(net135),
    .A2(_3162_),
    .B1(_3164_),
    .B2(_3153_),
    .C1(net207),
    .X(_0345_));
 sky130_fd_sc_hd__a21o_1 _6930_ (.A1(_2546_),
    .A2(_2547_),
    .B1(net133),
    .X(_3165_));
 sky130_fd_sc_hd__and3b_1 _6931_ (.A_N(_2548_),
    .B(_3165_),
    .C(_3513_),
    .X(_3166_));
 sky130_fd_sc_hd__nand3b_1 _6932_ (.A_N(_2517_),
    .B(_2558_),
    .C(_2559_),
    .Y(_3167_));
 sky130_fd_sc_hd__and3_1 _6933_ (.A(net101),
    .B(_2560_),
    .C(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__xnor2_1 _6934_ (.A(_2517_),
    .B(_2574_),
    .Y(_3169_));
 sky130_fd_sc_hd__or2_1 _6935_ (.A(net132),
    .B(net164),
    .X(_3170_));
 sky130_fd_sc_hd__o211a_1 _6936_ (.A1(net135),
    .A2(net117),
    .B1(_3517_),
    .C1(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__a221o_1 _6937_ (.A1(net126),
    .A2(_3570_),
    .B1(_3149_),
    .B2(_3169_),
    .C1(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__o31a_1 _6938_ (.A1(_3166_),
    .A2(_3168_),
    .A3(_3172_),
    .B1(net100),
    .X(_3173_));
 sky130_fd_sc_hd__xnor2_1 _6939_ (.A(_2519_),
    .B(_3113_),
    .Y(_3174_));
 sky130_fd_sc_hd__nor2_1 _6940_ (.A(net222),
    .B(_3174_),
    .Y(_3175_));
 sky130_fd_sc_hd__a31o_1 _6941_ (.A1(_3109_),
    .A2(_3110_),
    .A3(_3131_),
    .B1(net119),
    .X(_3176_));
 sky130_fd_sc_hd__o221a_1 _6942_ (.A1(net161),
    .A2(_2517_),
    .B1(_3175_),
    .B2(_3176_),
    .C1(_0502_),
    .X(_3177_));
 sky130_fd_sc_hd__o21ai_1 _6943_ (.A1(_3438_),
    .A2(net108),
    .B1(_2098_),
    .Y(_3178_));
 sky130_fd_sc_hd__a32o_1 _6944_ (.A1(net101),
    .A2(_2100_),
    .A3(_3178_),
    .B1(_3073_),
    .B2(net97),
    .X(_3179_));
 sky130_fd_sc_hd__nand2_1 _6945_ (.A(_2517_),
    .B(_2518_),
    .Y(_3180_));
 sky130_fd_sc_hd__nor2_1 _6946_ (.A(_0500_),
    .B(_2092_),
    .Y(_3181_));
 sky130_fd_sc_hd__a31o_1 _6947_ (.A1(_3513_),
    .A2(_2520_),
    .A3(_3180_),
    .B1(_3181_),
    .X(_3182_));
 sky130_fd_sc_hd__nand2b_1 _6948_ (.A_N(_2517_),
    .B(_2558_),
    .Y(_3183_));
 sky130_fd_sc_hd__xnor2_1 _6949_ (.A(_2517_),
    .B(_2536_),
    .Y(_3184_));
 sky130_fd_sc_hd__a32o_1 _6950_ (.A1(net101),
    .A2(_2592_),
    .A3(_3183_),
    .B1(_3184_),
    .B2(net97),
    .X(_3185_));
 sky130_fd_sc_hd__mux2_1 _6951_ (.A0(_3179_),
    .A1(_3185_),
    .S(net119),
    .X(_3186_));
 sky130_fd_sc_hd__or4_1 _6952_ (.A(_0585_),
    .B(_3171_),
    .C(_3182_),
    .D(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__o32a_1 _6953_ (.A1(net133),
    .A2(net828),
    .A3(_0586_),
    .B1(_3177_),
    .B2(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__a221o_1 _6954_ (.A1(_0428_),
    .A2(_0574_),
    .B1(_0578_),
    .B2(_3616_),
    .C1(net99),
    .X(_3189_));
 sky130_fd_sc_hd__o21ba_1 _6955_ (.A1(_0535_),
    .A2(_3188_),
    .B1_N(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__o21a_1 _6956_ (.A1(_3173_),
    .A2(_3190_),
    .B1(net105),
    .X(_3191_));
 sky130_fd_sc_hd__a21o_1 _6957_ (.A1(net32),
    .A2(net102),
    .B1(_3163_),
    .X(_3192_));
 sky130_fd_sc_hd__o221a_1 _6958_ (.A1(net133),
    .A2(_3162_),
    .B1(_3191_),
    .B2(_3192_),
    .C1(net208),
    .X(_0346_));
 sky130_fd_sc_hd__xnor2_1 _6959_ (.A(_2513_),
    .B(_2549_),
    .Y(_3193_));
 sky130_fd_sc_hd__nand2_1 _6960_ (.A(net101),
    .B(_2561_),
    .Y(_3194_));
 sky130_fd_sc_hd__a31o_1 _6961_ (.A1(_2092_),
    .A2(_2512_),
    .A3(_2560_),
    .B1(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__or2_1 _6962_ (.A(net130),
    .B(net164),
    .X(_3196_));
 sky130_fd_sc_hd__o211a_1 _6963_ (.A1(net133),
    .A2(net117),
    .B1(_3517_),
    .C1(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__a21oi_1 _6964_ (.A1(net123),
    .A2(_3570_),
    .B1(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hd__a2bb2o_1 _6965_ (.A1_N(_2512_),
    .A2_N(_2575_),
    .B1(_2576_),
    .B2(_2511_),
    .X(_3199_));
 sky130_fd_sc_hd__o22a_1 _6966_ (.A1(_3514_),
    .A2(_3193_),
    .B1(_3199_),
    .B2(_3148_),
    .X(_3200_));
 sky130_fd_sc_hd__a31o_1 _6967_ (.A1(_3195_),
    .A2(_3198_),
    .A3(_3200_),
    .B1(_0513_),
    .X(_3201_));
 sky130_fd_sc_hd__xnor2_1 _6968_ (.A(_3107_),
    .B(_3114_),
    .Y(_3202_));
 sky130_fd_sc_hd__nor2_1 _6969_ (.A(net222),
    .B(_3202_),
    .Y(_3203_));
 sky130_fd_sc_hd__a211o_1 _6970_ (.A1(_3103_),
    .A2(net222),
    .B1(_3203_),
    .C1(net119),
    .X(_3204_));
 sky130_fd_sc_hd__o211a_1 _6971_ (.A1(net161),
    .A2(_2513_),
    .B1(_3204_),
    .C1(_0502_),
    .X(_3205_));
 sky130_fd_sc_hd__or2_1 _6972_ (.A(_2099_),
    .B(_2101_),
    .X(_3206_));
 sky130_fd_sc_hd__a32o_1 _6973_ (.A1(net101),
    .A2(_2102_),
    .A3(_3206_),
    .B1(net243),
    .B2(net97),
    .X(_3207_));
 sky130_fd_sc_hd__and3_1 _6974_ (.A(_2513_),
    .B(_2514_),
    .C(_2520_),
    .X(_3208_));
 sky130_fd_sc_hd__o32a_1 _6975_ (.A1(_3514_),
    .A2(_2521_),
    .A3(_3208_),
    .B1(_0500_),
    .B2(_2036_),
    .X(_3209_));
 sky130_fd_sc_hd__a21oi_1 _6976_ (.A1(_2514_),
    .A2(_2536_),
    .B1(_2515_),
    .Y(_3210_));
 sky130_fd_sc_hd__xnor2_1 _6977_ (.A(_2512_),
    .B(_3210_),
    .Y(_3211_));
 sky130_fd_sc_hd__nand3_1 _6978_ (.A(_2092_),
    .B(_2512_),
    .C(_2592_),
    .Y(_3212_));
 sky130_fd_sc_hd__a32o_1 _6979_ (.A1(net101),
    .A2(_2593_),
    .A3(_3212_),
    .B1(_3211_),
    .B2(net97),
    .X(_3213_));
 sky130_fd_sc_hd__mux2_1 _6980_ (.A0(_3207_),
    .A1(_3213_),
    .S(net119),
    .X(_3214_));
 sky130_fd_sc_hd__or4b_1 _6981_ (.A(_0585_),
    .B(_3214_),
    .C(_3197_),
    .D_N(_3209_),
    .X(_3215_));
 sky130_fd_sc_hd__o32a_1 _6982_ (.A1(net132),
    .A2(net154),
    .A3(_0586_),
    .B1(_3205_),
    .B2(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__a221o_1 _6983_ (.A1(_0412_),
    .A2(_0574_),
    .B1(_0578_),
    .B2(_0462_),
    .C1(net99),
    .X(_3217_));
 sky130_fd_sc_hd__o21bai_1 _6984_ (.A1(_0535_),
    .A2(_3216_),
    .B1_N(_3217_),
    .Y(_3218_));
 sky130_fd_sc_hd__a21oi_1 _6985_ (.A1(_3201_),
    .A2(_3218_),
    .B1(net103),
    .Y(_3219_));
 sky130_fd_sc_hd__a21o_1 _6986_ (.A1(net33),
    .A2(net102),
    .B1(_3163_),
    .X(_3220_));
 sky130_fd_sc_hd__o221a_1 _6987_ (.A1(net132),
    .A2(_3162_),
    .B1(_3219_),
    .B2(_3220_),
    .C1(net208),
    .X(_0347_));
 sky130_fd_sc_hd__xnor2_1 _6988_ (.A(_2538_),
    .B(_2550_),
    .Y(_3221_));
 sky130_fd_sc_hd__nand2_1 _6989_ (.A(net101),
    .B(_2562_),
    .Y(_3222_));
 sky130_fd_sc_hd__a31o_1 _6990_ (.A1(_2036_),
    .A2(_2537_),
    .A3(_2561_),
    .B1(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__mux2_1 _6991_ (.A0(net127),
    .A1(net132),
    .S(\as1802.cond_inv ),
    .X(_3224_));
 sky130_fd_sc_hd__a22oi_1 _6992_ (.A1(net120),
    .A2(_3570_),
    .B1(_3224_),
    .B2(_3517_),
    .Y(_3225_));
 sky130_fd_sc_hd__nor2_1 _6993_ (.A(_2537_),
    .B(_2577_),
    .Y(_3226_));
 sky130_fd_sc_hd__a21o_1 _6994_ (.A1(_2537_),
    .A2(_2577_),
    .B1(_3148_),
    .X(_3227_));
 sky130_fd_sc_hd__o22a_1 _6995_ (.A1(_3514_),
    .A2(_3221_),
    .B1(_3226_),
    .B2(_3227_),
    .X(_3228_));
 sky130_fd_sc_hd__a31o_1 _6996_ (.A1(_3223_),
    .A2(_3225_),
    .A3(_3228_),
    .B1(_0513_),
    .X(_3229_));
 sky130_fd_sc_hd__o21ai_1 _6997_ (.A1(_3107_),
    .A2(_3114_),
    .B1(_3104_),
    .Y(_3230_));
 sky130_fd_sc_hd__xnor2_1 _6998_ (.A(_3116_),
    .B(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__nor2_1 _6999_ (.A(net222),
    .B(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__a21o_1 _7000_ (.A1(_3099_),
    .A2(net222),
    .B1(net119),
    .X(_3233_));
 sky130_fd_sc_hd__o221a_1 _7001_ (.A1(net162),
    .A2(_2538_),
    .B1(_3232_),
    .B2(_3233_),
    .C1(_0502_),
    .X(_3234_));
 sky130_fd_sc_hd__nand2_1 _7002_ (.A(_2102_),
    .B(_2103_),
    .Y(_3235_));
 sky130_fd_sc_hd__a32o_1 _7003_ (.A1(net101),
    .A2(_2104_),
    .A3(_3235_),
    .B1(net225),
    .B2(net98),
    .X(_3236_));
 sky130_fd_sc_hd__o21ai_1 _7004_ (.A1(_2522_),
    .A2(_2537_),
    .B1(_3513_),
    .Y(_3237_));
 sky130_fd_sc_hd__a21oi_1 _7005_ (.A1(_2522_),
    .A2(_2537_),
    .B1(_3237_),
    .Y(_3238_));
 sky130_fd_sc_hd__a2bb2o_1 _7006_ (.A1_N(_0500_),
    .A2_N(_1947_),
    .B1(_3224_),
    .B2(_3517_),
    .X(_3239_));
 sky130_fd_sc_hd__a21oi_1 _7007_ (.A1(_2511_),
    .A2(_3210_),
    .B1(_2509_),
    .Y(_3240_));
 sky130_fd_sc_hd__xor2_1 _7008_ (.A(_2537_),
    .B(_3240_),
    .X(_3241_));
 sky130_fd_sc_hd__nand3_1 _7009_ (.A(_2036_),
    .B(_2537_),
    .C(_2593_),
    .Y(_3242_));
 sky130_fd_sc_hd__a32o_1 _7010_ (.A1(net101),
    .A2(_2594_),
    .A3(_3242_),
    .B1(_3241_),
    .B2(net97),
    .X(_3243_));
 sky130_fd_sc_hd__mux2_1 _7011_ (.A0(_3236_),
    .A1(_3243_),
    .S(net119),
    .X(_3244_));
 sky130_fd_sc_hd__or4_1 _7012_ (.A(_0585_),
    .B(_3238_),
    .C(_3239_),
    .D(_3244_),
    .X(_3245_));
 sky130_fd_sc_hd__o32a_1 _7013_ (.A1(net130),
    .A2(net151),
    .A3(_0586_),
    .B1(_3234_),
    .B2(_3245_),
    .X(_3246_));
 sky130_fd_sc_hd__a221o_1 _7014_ (.A1(_0404_),
    .A2(_0574_),
    .B1(_0578_),
    .B2(_0472_),
    .C1(net99),
    .X(_3247_));
 sky130_fd_sc_hd__o21bai_1 _7015_ (.A1(_0535_),
    .A2(_3246_),
    .B1_N(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__a21oi_1 _7016_ (.A1(_3229_),
    .A2(_3248_),
    .B1(net103),
    .Y(_3249_));
 sky130_fd_sc_hd__a21o_1 _7017_ (.A1(net34),
    .A2(net102),
    .B1(_3163_),
    .X(_3250_));
 sky130_fd_sc_hd__o221a_1 _7018_ (.A1(net130),
    .A2(_3162_),
    .B1(_3249_),
    .B2(_3250_),
    .C1(net208),
    .X(_0348_));
 sky130_fd_sc_hd__nand2_1 _7019_ (.A(_2505_),
    .B(_2551_),
    .Y(_3251_));
 sky130_fd_sc_hd__and3_1 _7020_ (.A(_3513_),
    .B(_2552_),
    .C(_3251_),
    .X(_3252_));
 sky130_fd_sc_hd__or2_1 _7021_ (.A(_2504_),
    .B(_2578_),
    .X(_3253_));
 sky130_fd_sc_hd__nand2_1 _7022_ (.A(_2504_),
    .B(_2578_),
    .Y(_3254_));
 sky130_fd_sc_hd__and3_1 _7023_ (.A(_3149_),
    .B(_3253_),
    .C(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__a31o_1 _7024_ (.A1(_1947_),
    .A2(_2504_),
    .A3(_2562_),
    .B1(_3504_),
    .X(_3256_));
 sky130_fd_sc_hd__or2_1 _7025_ (.A(net126),
    .B(net164),
    .X(_3257_));
 sky130_fd_sc_hd__o211a_1 _7026_ (.A1(net130),
    .A2(net117),
    .B1(_3517_),
    .C1(_3257_),
    .X(_3258_));
 sky130_fd_sc_hd__a2bb2o_1 _7027_ (.A1_N(_2563_),
    .A2_N(_3256_),
    .B1(net135),
    .B2(_3570_),
    .X(_3259_));
 sky130_fd_sc_hd__o41a_1 _7028_ (.A1(_3252_),
    .A2(_3255_),
    .A3(_3258_),
    .A4(_3259_),
    .B1(net100),
    .X(_3260_));
 sky130_fd_sc_hd__and2_1 _7029_ (.A(_3091_),
    .B(_3131_),
    .X(_3261_));
 sky130_fd_sc_hd__xnor2_1 _7030_ (.A(_3094_),
    .B(_3117_),
    .Y(_3262_));
 sky130_fd_sc_hd__o21ai_1 _7031_ (.A1(net222),
    .A2(_3262_),
    .B1(net162),
    .Y(_3263_));
 sky130_fd_sc_hd__o221a_1 _7032_ (.A1(net162),
    .A2(_2505_),
    .B1(_3261_),
    .B2(_3263_),
    .C1(_0502_),
    .X(_3264_));
 sky130_fd_sc_hd__xnor2_1 _7033_ (.A(_2089_),
    .B(_2105_),
    .Y(_3265_));
 sky130_fd_sc_hd__a22o_1 _7034_ (.A1(net98),
    .A2(_2896_),
    .B1(_3265_),
    .B2(net101),
    .X(_3266_));
 sky130_fd_sc_hd__or3b_1 _7035_ (.A(_2504_),
    .B(_2507_),
    .C_N(_2523_),
    .X(_3267_));
 sky130_fd_sc_hd__a32o_1 _7036_ (.A1(_3513_),
    .A2(_2524_),
    .A3(_3267_),
    .B1(_0499_),
    .B2(_2005_),
    .X(_3268_));
 sky130_fd_sc_hd__a21o_1 _7037_ (.A1(_2506_),
    .A2(_3240_),
    .B1(_2508_),
    .X(_3269_));
 sky130_fd_sc_hd__or2_1 _7038_ (.A(_2504_),
    .B(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__nand2_1 _7039_ (.A(_2504_),
    .B(_3269_),
    .Y(_3271_));
 sky130_fd_sc_hd__and3_1 _7040_ (.A(_1947_),
    .B(_2504_),
    .C(_2594_),
    .X(_3272_));
 sky130_fd_sc_hd__nor2_1 _7041_ (.A(_2595_),
    .B(_3272_),
    .Y(_3273_));
 sky130_fd_sc_hd__a32o_1 _7042_ (.A1(net97),
    .A2(_3270_),
    .A3(_3271_),
    .B1(_3273_),
    .B2(net101),
    .X(_3274_));
 sky130_fd_sc_hd__mux2_1 _7043_ (.A0(_3266_),
    .A1(_3274_),
    .S(net119),
    .X(_3275_));
 sky130_fd_sc_hd__or4_1 _7044_ (.A(_0585_),
    .B(_3258_),
    .C(_3268_),
    .D(_3275_),
    .X(_3276_));
 sky130_fd_sc_hd__o32a_1 _7045_ (.A1(net127),
    .A2(net148),
    .A3(_0586_),
    .B1(_3264_),
    .B2(_3276_),
    .X(_3277_));
 sky130_fd_sc_hd__a221o_1 _7046_ (.A1(_0396_),
    .A2(_0574_),
    .B1(_0578_),
    .B2(_3608_),
    .C1(net99),
    .X(_3278_));
 sky130_fd_sc_hd__o21ba_1 _7047_ (.A1(_0535_),
    .A2(_3277_),
    .B1_N(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__o21a_1 _7048_ (.A1(_3260_),
    .A2(_3279_),
    .B1(net105),
    .X(_3280_));
 sky130_fd_sc_hd__a21o_1 _7049_ (.A1(net35),
    .A2(net102),
    .B1(_3163_),
    .X(_3281_));
 sky130_fd_sc_hd__o221a_1 _7050_ (.A1(net127),
    .A2(_3162_),
    .B1(_3280_),
    .B2(_3281_),
    .C1(net208),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _7051_ (.A(_2533_),
    .B(_2553_),
    .Y(_3282_));
 sky130_fd_sc_hd__o21a_1 _7052_ (.A1(_2533_),
    .A2(_2553_),
    .B1(_3513_),
    .X(_3283_));
 sky130_fd_sc_hd__o21ai_1 _7053_ (.A1(_2533_),
    .A2(_2564_),
    .B1(net101),
    .Y(_3284_));
 sky130_fd_sc_hd__a21o_1 _7054_ (.A1(_2533_),
    .A2(_2564_),
    .B1(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__a311o_1 _7055_ (.A1(_2503_),
    .A2(_2532_),
    .A3(_3254_),
    .B1(_3148_),
    .C1(_2579_),
    .X(_3286_));
 sky130_fd_sc_hd__or2_1 _7056_ (.A(net123),
    .B(net164),
    .X(_3287_));
 sky130_fd_sc_hd__o211a_1 _7057_ (.A1(net127),
    .A2(net117),
    .B1(_3517_),
    .C1(_3287_),
    .X(_3288_));
 sky130_fd_sc_hd__a221oi_1 _7058_ (.A1(net133),
    .A2(_3570_),
    .B1(_3282_),
    .B2(_3283_),
    .C1(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__a31o_1 _7059_ (.A1(_3285_),
    .A2(_3286_),
    .A3(_3289_),
    .B1(_0513_),
    .X(_3290_));
 sky130_fd_sc_hd__and2b_1 _7060_ (.A_N(_3086_),
    .B(_3131_),
    .X(_3291_));
 sky130_fd_sc_hd__a21oi_1 _7061_ (.A1(_3094_),
    .A2(_3117_),
    .B1(_3092_),
    .Y(_3292_));
 sky130_fd_sc_hd__xor2_1 _7062_ (.A(_3120_),
    .B(_3292_),
    .X(_3293_));
 sky130_fd_sc_hd__o21ai_1 _7063_ (.A1(_3131_),
    .A2(_3293_),
    .B1(net162),
    .Y(_3294_));
 sky130_fd_sc_hd__o221a_1 _7064_ (.A1(net162),
    .A2(_2532_),
    .B1(_3291_),
    .B2(_3294_),
    .C1(_0502_),
    .X(_3295_));
 sky130_fd_sc_hd__a21o_1 _7065_ (.A1(_2503_),
    .A2(_3271_),
    .B1(_2532_),
    .X(_3296_));
 sky130_fd_sc_hd__or3b_1 _7066_ (.A(_2502_),
    .B(_2533_),
    .C_N(_3271_),
    .X(_3297_));
 sky130_fd_sc_hd__a21o_1 _7067_ (.A1(_3296_),
    .A2(_3297_),
    .B1(net162),
    .X(_3298_));
 sky130_fd_sc_hd__o211a_1 _7068_ (.A1(_3439_),
    .A2(net227),
    .B1(_3298_),
    .C1(net98),
    .X(_3299_));
 sky130_fd_sc_hd__and3_1 _7069_ (.A(_2078_),
    .B(_2087_),
    .C(_2106_),
    .X(_3300_));
 sky130_fd_sc_hd__nor2_1 _7070_ (.A(_0500_),
    .B(_2166_),
    .Y(_3301_));
 sky130_fd_sc_hd__or2_1 _7071_ (.A(_2525_),
    .B(_2533_),
    .X(_3302_));
 sky130_fd_sc_hd__nand2_1 _7072_ (.A(_2525_),
    .B(_2533_),
    .Y(_3303_));
 sky130_fd_sc_hd__nor2_1 _7073_ (.A(_2107_),
    .B(_3300_),
    .Y(_3304_));
 sky130_fd_sc_hd__and2_1 _7074_ (.A(_2532_),
    .B(_2596_),
    .X(_3305_));
 sky130_fd_sc_hd__o21ai_1 _7075_ (.A1(_2532_),
    .A2(_2596_),
    .B1(net119),
    .Y(_3306_));
 sky130_fd_sc_hd__o221a_1 _7076_ (.A1(net119),
    .A2(_3304_),
    .B1(_3305_),
    .B2(_3306_),
    .C1(_3503_),
    .X(_3307_));
 sky130_fd_sc_hd__a311o_1 _7077_ (.A1(_3513_),
    .A2(_3302_),
    .A3(_3303_),
    .B1(_3307_),
    .C1(_3299_),
    .X(_3308_));
 sky130_fd_sc_hd__or4_1 _7078_ (.A(_0585_),
    .B(_3288_),
    .C(_3301_),
    .D(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__a2bb2o_1 _7079_ (.A1_N(_3295_),
    .A2_N(_3309_),
    .B1(_0585_),
    .B2(_2530_),
    .X(_3310_));
 sky130_fd_sc_hd__a221o_1 _7080_ (.A1(_0388_),
    .A2(_0574_),
    .B1(_0578_),
    .B2(_3600_),
    .C1(net100),
    .X(_3311_));
 sky130_fd_sc_hd__a21o_1 _7081_ (.A1(_0536_),
    .A2(_3310_),
    .B1(_3311_),
    .X(_3312_));
 sky130_fd_sc_hd__a21oi_1 _7082_ (.A1(_3290_),
    .A2(_3312_),
    .B1(net103),
    .Y(_3313_));
 sky130_fd_sc_hd__a21o_1 _7083_ (.A1(net36),
    .A2(net102),
    .B1(_3163_),
    .X(_3314_));
 sky130_fd_sc_hd__o221a_1 _7084_ (.A1(net126),
    .A2(_3162_),
    .B1(_3313_),
    .B2(_3314_),
    .C1(net208),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _7085_ (.A(_3082_),
    .B(_3122_),
    .Y(_3315_));
 sky130_fd_sc_hd__a21oi_1 _7086_ (.A1(_3123_),
    .A2(_3315_),
    .B1(net222),
    .Y(_3316_));
 sky130_fd_sc_hd__o311a_1 _7087_ (.A1(_3076_),
    .A2(_3082_),
    .A3(_3122_),
    .B1(_3129_),
    .C1(_3078_),
    .X(_3317_));
 sky130_fd_sc_hd__o21ai_1 _7088_ (.A1(_3316_),
    .A2(_3317_),
    .B1(net162),
    .Y(_3318_));
 sky130_fd_sc_hd__o211a_1 _7089_ (.A1(net162),
    .A2(_2535_),
    .B1(_3318_),
    .C1(_0502_),
    .X(_3319_));
 sky130_fd_sc_hd__or2_1 _7090_ (.A(_3439_),
    .B(_2777_),
    .X(_3320_));
 sky130_fd_sc_hd__a21o_1 _7091_ (.A1(_2500_),
    .A2(_3296_),
    .B1(_2535_),
    .X(_3321_));
 sky130_fd_sc_hd__or3b_1 _7092_ (.A(_2499_),
    .B(_2534_),
    .C_N(_3296_),
    .X(_3322_));
 sky130_fd_sc_hd__a21o_1 _7093_ (.A1(_3321_),
    .A2(_3322_),
    .B1(net162),
    .X(_3323_));
 sky130_fd_sc_hd__a21oi_1 _7094_ (.A1(_2076_),
    .A2(_2108_),
    .B1(_2107_),
    .Y(_3324_));
 sky130_fd_sc_hd__or3b_1 _7095_ (.A(_3136_),
    .B(_3324_),
    .C_N(_2109_),
    .X(_3325_));
 sky130_fd_sc_hd__xnor2_1 _7096_ (.A(_2526_),
    .B(_2534_),
    .Y(_3326_));
 sky130_fd_sc_hd__mux2_1 _7097_ (.A0(net120),
    .A1(net126),
    .S(\as1802.cond_inv ),
    .X(_3327_));
 sky130_fd_sc_hd__nand2_1 _7098_ (.A(_3517_),
    .B(_3327_),
    .Y(_3328_));
 sky130_fd_sc_hd__o221a_1 _7099_ (.A1(_0500_),
    .A2(_2222_),
    .B1(_3326_),
    .B2(_3514_),
    .C1(_0586_),
    .X(_3329_));
 sky130_fd_sc_hd__and3_1 _7100_ (.A(_2166_),
    .B(_2534_),
    .C(_2597_),
    .X(_3330_));
 sky130_fd_sc_hd__or3_1 _7101_ (.A(_3505_),
    .B(_2598_),
    .C(_3330_),
    .X(_3331_));
 sky130_fd_sc_hd__nand4_1 _7102_ (.A(_3325_),
    .B(_3328_),
    .C(_3329_),
    .D(_3331_),
    .Y(_3332_));
 sky130_fd_sc_hd__a31o_1 _7103_ (.A1(net97),
    .A2(_3320_),
    .A3(_3323_),
    .B1(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__o31a_1 _7104_ (.A1(net123),
    .A2(net142),
    .A3(_0586_),
    .B1(_0579_),
    .X(_3334_));
 sky130_fd_sc_hd__o21ai_1 _7105_ (.A1(_3319_),
    .A2(_3333_),
    .B1(_3334_),
    .Y(_3335_));
 sky130_fd_sc_hd__a21o_1 _7106_ (.A1(net163),
    .A2(_3592_),
    .B1(_0536_),
    .X(_3336_));
 sky130_fd_sc_hd__a221o_1 _7107_ (.A1(_0441_),
    .A2(_0574_),
    .B1(_3335_),
    .B2(_3336_),
    .C1(net100),
    .X(_3337_));
 sky130_fd_sc_hd__xnor2_1 _7108_ (.A(_2534_),
    .B(_2554_),
    .Y(_3338_));
 sky130_fd_sc_hd__and3_1 _7109_ (.A(_2166_),
    .B(_2534_),
    .C(_2565_),
    .X(_3339_));
 sky130_fd_sc_hd__xnor2_1 _7110_ (.A(_2535_),
    .B(_2580_),
    .Y(_3340_));
 sky130_fd_sc_hd__o32a_1 _7111_ (.A1(_3504_),
    .A2(_2566_),
    .A3(_3339_),
    .B1(_3571_),
    .B2(_3436_),
    .X(_3341_));
 sky130_fd_sc_hd__o22a_1 _7112_ (.A1(_3514_),
    .A2(_3338_),
    .B1(_3340_),
    .B2(_3148_),
    .X(_3342_));
 sky130_fd_sc_hd__a31o_1 _7113_ (.A1(_3328_),
    .A2(_3341_),
    .A3(_3342_),
    .B1(_0513_),
    .X(_3343_));
 sky130_fd_sc_hd__a21oi_1 _7114_ (.A1(_3337_),
    .A2(_3343_),
    .B1(net103),
    .Y(_3344_));
 sky130_fd_sc_hd__a21o_1 _7115_ (.A1(net37),
    .A2(net102),
    .B1(_3163_),
    .X(_3345_));
 sky130_fd_sc_hd__o221a_1 _7116_ (.A1(net123),
    .A2(_3162_),
    .B1(_3344_),
    .B2(_3345_),
    .C1(net208),
    .X(_0351_));
 sky130_fd_sc_hd__a21oi_1 _7117_ (.A1(_2494_),
    .A2(_2555_),
    .B1(_3514_),
    .Y(_3346_));
 sky130_fd_sc_hd__o21a_1 _7118_ (.A1(_2494_),
    .A2(_2555_),
    .B1(_3346_),
    .X(_3347_));
 sky130_fd_sc_hd__a21oi_1 _7119_ (.A1(_2494_),
    .A2(_2567_),
    .B1(_3504_),
    .Y(_3348_));
 sky130_fd_sc_hd__o21a_1 _7120_ (.A1(_2494_),
    .A2(_2567_),
    .B1(_3348_),
    .X(_3349_));
 sky130_fd_sc_hd__nor2_1 _7121_ (.A(_2494_),
    .B(_2581_),
    .Y(_3350_));
 sky130_fd_sc_hd__or2_1 _7122_ (.A(_2582_),
    .B(_3350_),
    .X(_3351_));
 sky130_fd_sc_hd__and3_1 _7123_ (.A(net123),
    .B(_3515_),
    .C(_3563_),
    .X(_3352_));
 sky130_fd_sc_hd__a21o_1 _7124_ (.A1(net130),
    .A2(_3570_),
    .B1(_3352_),
    .X(_3353_));
 sky130_fd_sc_hd__a31o_1 _7125_ (.A1(net871),
    .A2(net117),
    .A3(_3517_),
    .B1(_3353_),
    .X(_3354_));
 sky130_fd_sc_hd__a21o_1 _7126_ (.A1(_3149_),
    .A2(_3351_),
    .B1(_3354_),
    .X(_3355_));
 sky130_fd_sc_hd__o31a_1 _7127_ (.A1(_3347_),
    .A2(_3349_),
    .A3(_3355_),
    .B1(net100),
    .X(_3356_));
 sky130_fd_sc_hd__a21oi_1 _7128_ (.A1(_3081_),
    .A2(_3121_),
    .B1(_3079_),
    .Y(_3357_));
 sky130_fd_sc_hd__xnor2_1 _7129_ (.A(_3076_),
    .B(_3357_),
    .Y(_3358_));
 sky130_fd_sc_hd__nor2_1 _7130_ (.A(_3131_),
    .B(_3358_),
    .Y(_3359_));
 sky130_fd_sc_hd__a21o_1 _7131_ (.A1(_3075_),
    .A2(_3131_),
    .B1(net119),
    .X(_3360_));
 sky130_fd_sc_hd__o221a_1 _7132_ (.A1(net162),
    .A2(_2495_),
    .B1(_3359_),
    .B2(_3360_),
    .C1(_0502_),
    .X(_3361_));
 sky130_fd_sc_hd__a21oi_1 _7133_ (.A1(_2497_),
    .A2(_3321_),
    .B1(_2494_),
    .Y(_3362_));
 sky130_fd_sc_hd__a31o_1 _7134_ (.A1(_2494_),
    .A2(_2497_),
    .A3(_3321_),
    .B1(net57),
    .X(_3363_));
 sky130_fd_sc_hd__o221a_1 _7135_ (.A1(net119),
    .A2(_2715_),
    .B1(_3362_),
    .B2(_3363_),
    .C1(net97),
    .X(_3364_));
 sky130_fd_sc_hd__o211a_1 _7136_ (.A1(_2057_),
    .A2(_2058_),
    .B1(_2076_),
    .C1(_2109_),
    .X(_3365_));
 sky130_fd_sc_hd__or2_1 _7137_ (.A(_2494_),
    .B(_2527_),
    .X(_3366_));
 sky130_fd_sc_hd__a311o_1 _7138_ (.A1(net120),
    .A2(net139),
    .A3(_0499_),
    .B1(_0585_),
    .C1(_3352_),
    .X(_3367_));
 sky130_fd_sc_hd__a31o_1 _7139_ (.A1(_3513_),
    .A2(_2528_),
    .A3(_3366_),
    .B1(_3367_),
    .X(_3368_));
 sky130_fd_sc_hd__o21ai_1 _7140_ (.A1(_2110_),
    .A2(_3365_),
    .B1(net57),
    .Y(_3369_));
 sky130_fd_sc_hd__o21ai_1 _7141_ (.A1(_2495_),
    .A2(_2599_),
    .B1(net119),
    .Y(_3370_));
 sky130_fd_sc_hd__a21o_1 _7142_ (.A1(_2495_),
    .A2(_2599_),
    .B1(_3370_),
    .X(_3371_));
 sky130_fd_sc_hd__a311o_1 _7143_ (.A1(net101),
    .A2(_3369_),
    .A3(_3371_),
    .B1(_3364_),
    .C1(_3368_),
    .X(_3372_));
 sky130_fd_sc_hd__a2bb2o_1 _7144_ (.A1_N(_3361_),
    .A2_N(_3372_),
    .B1(_0585_),
    .B2(_2492_),
    .X(_3373_));
 sky130_fd_sc_hd__a221o_1 _7145_ (.A1(_0451_),
    .A2(_0574_),
    .B1(_0578_),
    .B2(_0485_),
    .C1(net100),
    .X(_3374_));
 sky130_fd_sc_hd__a21oi_1 _7146_ (.A1(_0536_),
    .A2(_3373_),
    .B1(_3374_),
    .Y(_3375_));
 sky130_fd_sc_hd__o21a_1 _7147_ (.A1(_3356_),
    .A2(_3375_),
    .B1(net105),
    .X(_3376_));
 sky130_fd_sc_hd__a21o_1 _7148_ (.A1(net38),
    .A2(net103),
    .B1(_3163_),
    .X(_3377_));
 sky130_fd_sc_hd__o221a_1 _7149_ (.A1(net120),
    .A2(_3162_),
    .B1(_3376_),
    .B2(_3377_),
    .C1(net208),
    .X(_0352_));
 sky130_fd_sc_hd__and3_4 _7150_ (.A(_0635_),
    .B(_1256_),
    .C(_1316_),
    .X(_3378_));
 sky130_fd_sc_hd__and3_4 _7151_ (.A(_0704_),
    .B(_1259_),
    .C(_1318_),
    .X(_3379_));
 sky130_fd_sc_hd__mux2_1 _7152_ (.A0(net672),
    .A1(_0926_),
    .S(_3379_),
    .X(_3380_));
 sky130_fd_sc_hd__mux2_1 _7153_ (.A0(net673),
    .A1(_0652_),
    .S(_3378_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _7154_ (.A0(net676),
    .A1(_0974_),
    .S(_3379_),
    .X(_3381_));
 sky130_fd_sc_hd__mux2_1 _7155_ (.A0(_3381_),
    .A1(_0934_),
    .S(_3378_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _7156_ (.A0(net529),
    .A1(_1022_),
    .S(_3379_),
    .X(_3382_));
 sky130_fd_sc_hd__mux2_1 _7157_ (.A0(net530),
    .A1(_0982_),
    .S(_3378_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _7158_ (.A0(net448),
    .A1(_1067_),
    .S(_3379_),
    .X(_3383_));
 sky130_fd_sc_hd__mux2_1 _7159_ (.A0(net449),
    .A1(_1030_),
    .S(_3378_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _7160_ (.A0(net463),
    .A1(_1117_),
    .S(_3379_),
    .X(_3384_));
 sky130_fd_sc_hd__mux2_1 _7161_ (.A0(_3384_),
    .A1(_1075_),
    .S(_3378_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _7162_ (.A0(net684),
    .A1(_1165_),
    .S(_3379_),
    .X(_3385_));
 sky130_fd_sc_hd__mux2_1 _7163_ (.A0(net685),
    .A1(_1125_),
    .S(_3378_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _7164_ (.A0(net460),
    .A1(_1214_),
    .S(_3379_),
    .X(_3386_));
 sky130_fd_sc_hd__mux2_1 _7165_ (.A0(_3386_),
    .A1(_1172_),
    .S(_3378_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _7166_ (.A0(net419),
    .A1(_1253_),
    .S(_3379_),
    .X(_3387_));
 sky130_fd_sc_hd__mux2_1 _7167_ (.A0(_3387_),
    .A1(_1219_),
    .S(_3378_),
    .X(_0360_));
 sky130_fd_sc_hd__or4b_1 _7168_ (.A(_0575_),
    .B(_2316_),
    .C(_2657_),
    .D_N(_2654_),
    .X(_3388_));
 sky130_fd_sc_hd__or3_1 _7169_ (.A(_2279_),
    .B(_2282_),
    .C(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__nand3b_1 _7170_ (.A_N(_2284_),
    .B(_2315_),
    .C(_2317_),
    .Y(_3390_));
 sky130_fd_sc_hd__or3_1 _7171_ (.A(_2313_),
    .B(_3389_),
    .C(_3390_),
    .X(_3391_));
 sky130_fd_sc_hd__o2bb2a_1 _7172_ (.A1_N(net100),
    .A2_N(_2624_),
    .B1(net164),
    .B2(_3525_),
    .X(_3392_));
 sky130_fd_sc_hd__a21oi_1 _7173_ (.A1(_3524_),
    .A2(_3392_),
    .B1(net172),
    .Y(_3393_));
 sky130_fd_sc_hd__mux2_1 _7174_ (.A0(_3393_),
    .A1(net366),
    .S(net825),
    .X(_0361_));
 sky130_fd_sc_hd__and3_4 _7175_ (.A(_0635_),
    .B(_1257_),
    .C(_1270_),
    .X(_3394_));
 sky130_fd_sc_hd__and3_4 _7176_ (.A(_0704_),
    .B(_1260_),
    .C(_1273_),
    .X(_3395_));
 sky130_fd_sc_hd__mux2_1 _7177_ (.A0(net840),
    .A1(_0926_),
    .S(_3395_),
    .X(_3396_));
 sky130_fd_sc_hd__mux2_1 _7178_ (.A0(_3396_),
    .A1(_0652_),
    .S(_3394_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _7179_ (.A0(net867),
    .A1(_0974_),
    .S(_3395_),
    .X(_3397_));
 sky130_fd_sc_hd__mux2_1 _7180_ (.A0(_3397_),
    .A1(_0934_),
    .S(_3394_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _7181_ (.A0(net874),
    .A1(_1022_),
    .S(_3395_),
    .X(_3398_));
 sky130_fd_sc_hd__mux2_1 _7182_ (.A0(_3398_),
    .A1(_0982_),
    .S(_3394_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _7183_ (.A0(net844),
    .A1(_1067_),
    .S(_3395_),
    .X(_3399_));
 sky130_fd_sc_hd__mux2_1 _7184_ (.A0(net845),
    .A1(_1030_),
    .S(_3394_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _7185_ (.A0(net868),
    .A1(_1117_),
    .S(_3395_),
    .X(_3400_));
 sky130_fd_sc_hd__mux2_1 _7186_ (.A0(_3400_),
    .A1(_1075_),
    .S(_3394_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _7187_ (.A0(net838),
    .A1(_1165_),
    .S(_3395_),
    .X(_3401_));
 sky130_fd_sc_hd__mux2_1 _7188_ (.A0(_3401_),
    .A1(_1125_),
    .S(_3394_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _7189_ (.A0(net869),
    .A1(_1214_),
    .S(_3395_),
    .X(_3402_));
 sky130_fd_sc_hd__mux2_1 _7190_ (.A0(_3402_),
    .A1(_1172_),
    .S(_3394_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _7191_ (.A0(net863),
    .A1(_1253_),
    .S(_3395_),
    .X(_3403_));
 sky130_fd_sc_hd__mux2_1 _7192_ (.A0(_3403_),
    .A1(_1219_),
    .S(_3394_),
    .X(_0369_));
 sky130_fd_sc_hd__and3_4 _7193_ (.A(_0635_),
    .B(_1270_),
    .C(_1316_),
    .X(_3404_));
 sky130_fd_sc_hd__and3_4 _7194_ (.A(_0704_),
    .B(_1273_),
    .C(_1318_),
    .X(_3405_));
 sky130_fd_sc_hd__mux2_1 _7195_ (.A0(net422),
    .A1(_0926_),
    .S(_3405_),
    .X(_3406_));
 sky130_fd_sc_hd__mux2_1 _7196_ (.A0(net423),
    .A1(_0652_),
    .S(_3404_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _7197_ (.A0(net418),
    .A1(_0974_),
    .S(_3405_),
    .X(_3407_));
 sky130_fd_sc_hd__mux2_1 _7198_ (.A0(_3407_),
    .A1(_0934_),
    .S(_3404_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _7199_ (.A0(net437),
    .A1(_1022_),
    .S(_3405_),
    .X(_3408_));
 sky130_fd_sc_hd__mux2_1 _7200_ (.A0(net438),
    .A1(_0982_),
    .S(_3404_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _7201_ (.A0(net454),
    .A1(_1067_),
    .S(_3405_),
    .X(_3409_));
 sky130_fd_sc_hd__mux2_1 _7202_ (.A0(net455),
    .A1(_1030_),
    .S(_3404_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _7203_ (.A0(net391),
    .A1(_1117_),
    .S(_3405_),
    .X(_3410_));
 sky130_fd_sc_hd__mux2_1 _7204_ (.A0(_3410_),
    .A1(_1075_),
    .S(_3404_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _7205_ (.A0(net568),
    .A1(_1165_),
    .S(_3405_),
    .X(_3411_));
 sky130_fd_sc_hd__mux2_1 _7206_ (.A0(net569),
    .A1(_1125_),
    .S(_3404_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _7207_ (.A0(net406),
    .A1(_1214_),
    .S(_3405_),
    .X(_3412_));
 sky130_fd_sc_hd__mux2_1 _7208_ (.A0(_3412_),
    .A1(_1172_),
    .S(_3404_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _7209_ (.A0(net524),
    .A1(_1253_),
    .S(_3405_),
    .X(_3413_));
 sky130_fd_sc_hd__mux2_1 _7210_ (.A0(_3413_),
    .A1(_1219_),
    .S(_3404_),
    .X(_0377_));
 sky130_fd_sc_hd__and3b_4 _7211_ (.A_N(_0633_),
    .B(_0635_),
    .C(_1270_),
    .X(_3414_));
 sky130_fd_sc_hd__and3_4 _7212_ (.A(_0702_),
    .B(_0704_),
    .C(_1273_),
    .X(_3415_));
 sky130_fd_sc_hd__mux2_1 _7213_ (.A0(net383),
    .A1(_0926_),
    .S(_3415_),
    .X(_3416_));
 sky130_fd_sc_hd__mux2_1 _7214_ (.A0(net384),
    .A1(_0652_),
    .S(_3414_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _7215_ (.A0(net598),
    .A1(_0974_),
    .S(_3415_),
    .X(_3417_));
 sky130_fd_sc_hd__mux2_1 _7216_ (.A0(_3417_),
    .A1(_0934_),
    .S(_3414_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _7217_ (.A0(net508),
    .A1(_1022_),
    .S(_3415_),
    .X(_3418_));
 sky130_fd_sc_hd__mux2_1 _7218_ (.A0(net509),
    .A1(_0982_),
    .S(_3414_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _7219_ (.A0(net584),
    .A1(_1067_),
    .S(_3415_),
    .X(_3419_));
 sky130_fd_sc_hd__mux2_1 _7220_ (.A0(net585),
    .A1(_1030_),
    .S(_3414_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _7221_ (.A0(net445),
    .A1(_1117_),
    .S(_3415_),
    .X(_3420_));
 sky130_fd_sc_hd__mux2_1 _7222_ (.A0(_3420_),
    .A1(_1075_),
    .S(_3414_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _7223_ (.A0(net396),
    .A1(_1165_),
    .S(_3415_),
    .X(_3421_));
 sky130_fd_sc_hd__mux2_1 _7224_ (.A0(net397),
    .A1(_1125_),
    .S(_3414_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _7225_ (.A0(net621),
    .A1(_1214_),
    .S(_3415_),
    .X(_3422_));
 sky130_fd_sc_hd__mux2_1 _7226_ (.A0(_3422_),
    .A1(_1172_),
    .S(_3414_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _7227_ (.A0(net484),
    .A1(_1253_),
    .S(_3415_),
    .X(_3423_));
 sky130_fd_sc_hd__mux2_1 _7228_ (.A0(_3423_),
    .A1(_1219_),
    .S(_3414_),
    .X(_0385_));
 sky130_fd_sc_hd__o2111a_1 _7229_ (.A1(net172),
    .A2(_3524_),
    .B1(_3539_),
    .C1(_0582_),
    .D1(net209),
    .X(_3424_));
 sky130_fd_sc_hd__or4_1 _7230_ (.A(net164),
    .B(_3525_),
    .C(_3580_),
    .D(_2621_),
    .X(_3425_));
 sky130_fd_sc_hd__and4_1 _7231_ (.A(_2317_),
    .B(_2610_),
    .C(_3424_),
    .D(_3425_),
    .X(_3426_));
 sky130_fd_sc_hd__and3_1 _7232_ (.A(_2280_),
    .B(_2314_),
    .C(_3426_),
    .X(_3427_));
 sky130_fd_sc_hd__or3b_1 _7233_ (.A(_2312_),
    .B(_3389_),
    .C_N(_3427_),
    .X(_3428_));
 sky130_fd_sc_hd__o21ai_1 _7234_ (.A1(\as1802.instr_latch[7] ),
    .A2(_3493_),
    .B1(_3525_),
    .Y(_3429_));
 sky130_fd_sc_hd__a31o_1 _7235_ (.A1(net95),
    .A2(_3580_),
    .A3(_0513_),
    .B1(_0526_),
    .X(_3430_));
 sky130_fd_sc_hd__o21a_1 _7236_ (.A1(_3429_),
    .A2(_3430_),
    .B1(net88),
    .X(_3431_));
 sky130_fd_sc_hd__mux2_1 _7237_ (.A0(_3431_),
    .A1(net276),
    .S(_3428_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _7238_ (.A0(_0598_),
    .A1(net431),
    .S(_0595_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _7239_ (.A0(net329),
    .A1(net278),
    .S(_0595_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _7240_ (.A0(net822),
    .A1(net819),
    .S(_0595_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _7241_ (.A0(_0609_),
    .A1(net472),
    .S(_0595_),
    .X(_0296_));
 sky130_fd_sc_hd__o211a_1 _7242_ (.A1(net31),
    .A2(_1567_),
    .B1(_1568_),
    .C1(net207),
    .X(_0310_));
 sky130_fd_sc_hd__o211a_1 _7243_ (.A1(net32),
    .A2(_1567_),
    .B1(_1569_),
    .C1(net207),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _7244_ (.A(net206),
    .B(_1570_),
    .X(_0312_));
 sky130_fd_sc_hd__o211a_1 _7245_ (.A1(net34),
    .A2(_1567_),
    .B1(_1571_),
    .C1(net208),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _7246_ (.A0(net317),
    .A1(net284),
    .S(_0613_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _7247_ (.A0(_0617_),
    .A1(net742),
    .S(_0613_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _7248_ (.A0(_0619_),
    .A1(net776),
    .S(_0613_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _7249_ (.A0(_0621_),
    .A1(net310),
    .S(_0613_),
    .X(_0333_));
 sky130_fd_sc_hd__dfxtp_1 _7250_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0028_),
    .Q(\as1802.regs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7251_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0029_),
    .Q(\as1802.regs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7252_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0030_),
    .Q(\as1802.regs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7253_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0031_),
    .Q(\as1802.regs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7254_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0032_),
    .Q(\as1802.regs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7255_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0033_),
    .Q(\as1802.regs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7256_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0034_),
    .Q(\as1802.regs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7257_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0035_),
    .Q(\as1802.regs[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _7258_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(net289),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_2 _7259_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(net818),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _7260_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0038_),
    .Q(\as1802.regs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7261_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0039_),
    .Q(\as1802.regs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7262_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0040_),
    .Q(\as1802.regs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7263_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0041_),
    .Q(\as1802.regs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7264_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0042_),
    .Q(\as1802.regs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7265_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0043_),
    .Q(\as1802.regs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7266_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0044_),
    .Q(\as1802.regs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7267_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0045_),
    .Q(\as1802.regs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7268_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0046_),
    .Q(\as1802.regs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7269_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0047_),
    .Q(\as1802.regs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7270_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0048_),
    .Q(\as1802.regs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7271_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0049_),
    .Q(\as1802.regs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7272_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0050_),
    .Q(\as1802.regs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7273_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0051_),
    .Q(\as1802.regs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7274_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0052_),
    .Q(\as1802.regs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7275_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0053_),
    .Q(\as1802.regs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7276_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0054_),
    .Q(\as1802.regs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7277_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0055_),
    .Q(\as1802.regs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7278_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0056_),
    .Q(\as1802.regs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7279_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0057_),
    .Q(\as1802.regs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7280_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0058_),
    .Q(\as1802.regs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7281_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0059_),
    .Q(\as1802.regs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7282_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0060_),
    .Q(\as1802.regs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7283_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0061_),
    .Q(\as1802.regs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7284_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0062_),
    .Q(\as1802.regs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7285_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0063_),
    .Q(\as1802.regs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7286_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0064_),
    .Q(\as1802.regs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7287_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0065_),
    .Q(\as1802.regs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7288_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0066_),
    .Q(\as1802.regs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7289_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0067_),
    .Q(\as1802.regs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7290_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0068_),
    .Q(\as1802.regs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7291_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0069_),
    .Q(\as1802.regs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7292_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0070_),
    .Q(\as1802.regs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7293_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0071_),
    .Q(\as1802.regs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7294_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0072_),
    .Q(\as1802.regs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7295_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0073_),
    .Q(\as1802.regs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7296_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0074_),
    .Q(\as1802.regs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7297_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0075_),
    .Q(\as1802.regs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7298_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0076_),
    .Q(\as1802.regs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7299_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0077_),
    .Q(\as1802.regs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7300_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0078_),
    .Q(\as1802.regs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7301_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0079_),
    .Q(\as1802.regs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7302_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0080_),
    .Q(\as1802.regs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7303_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0081_),
    .Q(\as1802.regs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7304_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0082_),
    .Q(\as1802.regs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7305_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0083_),
    .Q(\as1802.regs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7306_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0084_),
    .Q(\as1802.regs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7307_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0085_),
    .Q(\as1802.regs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7308_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0086_),
    .Q(\as1802.regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7309_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0087_),
    .Q(\as1802.regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7310_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0088_),
    .Q(\as1802.regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7311_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0089_),
    .Q(\as1802.regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7312_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0090_),
    .Q(\as1802.regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7313_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net772),
    .Q(\as1802.regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7314_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0092_),
    .Q(\as1802.regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7315_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0093_),
    .Q(\as1802.regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7316_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0094_),
    .Q(\as1802.regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7317_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0095_),
    .Q(\as1802.regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7318_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0096_),
    .Q(\as1802.regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7319_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0097_),
    .Q(\as1802.regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7320_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0098_),
    .Q(\as1802.regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7321_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net469),
    .Q(\as1802.regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7322_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0100_),
    .Q(\as1802.regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7323_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0101_),
    .Q(\as1802.regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7324_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0102_),
    .Q(\as1802.regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7325_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0103_),
    .Q(\as1802.regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7326_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net631),
    .Q(\as1802.regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7327_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0105_),
    .Q(\as1802.regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7328_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0106_),
    .Q(\as1802.regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7329_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net783),
    .Q(\as1802.regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7330_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0108_),
    .Q(\as1802.regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7331_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0109_),
    .Q(\as1802.regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7332_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0110_),
    .Q(\as1802.regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7333_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0111_),
    .Q(\as1802.regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7334_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0112_),
    .Q(\as1802.regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7335_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0113_),
    .Q(\as1802.regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7336_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0114_),
    .Q(\as1802.regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7337_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net382),
    .Q(\as1802.regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7338_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0116_),
    .Q(\as1802.regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7339_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0117_),
    .Q(\as1802.regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_4 _7340_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net432),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_4 _7341_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net279),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_2 _7342_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net820),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_2 _7343_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net535),
    .Q(_0007_));
 sky130_fd_sc_hd__dfxtp_2 _7344_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0118_),
    .Q(\as1802.regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7345_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0119_),
    .Q(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7346_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0120_),
    .Q(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _7347_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0121_),
    .Q(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7348_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0122_),
    .Q(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7349_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net848),
    .Q(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7350_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0124_),
    .Q(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _7351_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0125_),
    .Q(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7352_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0126_),
    .Q(\as1802.regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7353_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0127_),
    .Q(\as1802.regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7354_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0128_),
    .Q(\as1802.regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7355_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0129_),
    .Q(\as1802.regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7356_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0130_),
    .Q(\as1802.regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7357_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net760),
    .Q(\as1802.regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7358_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0132_),
    .Q(\as1802.regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7359_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0133_),
    .Q(\as1802.regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_4 _7360_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0134_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_4 _7361_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0135_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_4 _7362_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0136_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_4 _7363_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0137_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _7364_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0138_),
    .Q(\as1802.regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7365_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0139_),
    .Q(\as1802.regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7366_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net722),
    .Q(\as1802.regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7367_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0141_),
    .Q(\as1802.regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7368_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0142_),
    .Q(\as1802.regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7369_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net565),
    .Q(\as1802.regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7370_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net805),
    .Q(\as1802.regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7371_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0145_),
    .Q(\as1802.regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7372_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0146_),
    .Q(\as1802.regs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7373_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0147_),
    .Q(\as1802.regs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7374_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0148_),
    .Q(\as1802.regs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7375_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0149_),
    .Q(\as1802.regs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7376_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0150_),
    .Q(\as1802.regs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7377_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0151_),
    .Q(\as1802.regs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7378_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0152_),
    .Q(\as1802.regs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7379_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0153_),
    .Q(\as1802.regs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7380_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net751),
    .Q(\as1802.regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7381_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0155_),
    .Q(\as1802.regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7382_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net576),
    .Q(\as1802.regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7383_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0157_),
    .Q(\as1802.regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7384_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0158_),
    .Q(\as1802.regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7385_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net739),
    .Q(\as1802.regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7386_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0160_),
    .Q(\as1802.regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7387_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0161_),
    .Q(\as1802.regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7388_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net746),
    .Q(\as1802.regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7389_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0163_),
    .Q(\as1802.regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7390_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net477),
    .Q(\as1802.regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7391_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0165_),
    .Q(\as1802.regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7392_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0166_),
    .Q(\as1802.regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7393_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net634),
    .Q(\as1802.regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7394_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net808),
    .Q(\as1802.regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7395_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0169_),
    .Q(\as1802.regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7396_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0170_),
    .Q(\as1802.regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7397_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0171_),
    .Q(\as1802.regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7398_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net588),
    .Q(\as1802.regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7399_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0173_),
    .Q(\as1802.regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7400_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0174_),
    .Q(\as1802.regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7401_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net600),
    .Q(\as1802.regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7402_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0176_),
    .Q(\as1802.regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7403_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0177_),
    .Q(\as1802.regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7404_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0178_),
    .Q(\as1802.regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7405_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0179_),
    .Q(\as1802.regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7406_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net494),
    .Q(\as1802.regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7407_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0181_),
    .Q(\as1802.regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7408_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0182_),
    .Q(\as1802.regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7409_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net717),
    .Q(\as1802.regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7410_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net725),
    .Q(\as1802.regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7411_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0185_),
    .Q(\as1802.regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7412_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0186_),
    .Q(\as1802.regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7413_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0187_),
    .Q(\as1802.regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7414_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net554),
    .Q(\as1802.regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7415_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0189_),
    .Q(\as1802.regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7416_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0190_),
    .Q(\as1802.regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7417_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net609),
    .Q(\as1802.regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7418_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0192_),
    .Q(\as1802.regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7419_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0193_),
    .Q(\as1802.regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7420_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0194_),
    .Q(\as1802.regs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7421_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0195_),
    .Q(\as1802.regs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7422_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0196_),
    .Q(\as1802.regs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7423_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0197_),
    .Q(\as1802.regs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7424_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0198_),
    .Q(\as1802.regs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7425_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net623),
    .Q(\as1802.regs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7426_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0200_),
    .Q(\as1802.regs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7427_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0201_),
    .Q(\as1802.regs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7428_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0202_),
    .Q(\as1802.regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7429_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0203_),
    .Q(\as1802.regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7430_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net488),
    .Q(\as1802.regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7431_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0205_),
    .Q(\as1802.regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7432_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0206_),
    .Q(\as1802.regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7433_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net503),
    .Q(\as1802.regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7434_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0208_),
    .Q(\as1802.regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7435_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0209_),
    .Q(\as1802.regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7436_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net619),
    .Q(\as1802.regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7437_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0211_),
    .Q(\as1802.regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7438_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net458),
    .Q(\as1802.regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7439_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0213_),
    .Q(\as1802.regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7440_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0214_),
    .Q(\as1802.regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7441_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net638),
    .Q(\as1802.regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7442_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0216_),
    .Q(\as1802.regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7443_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0217_),
    .Q(\as1802.regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7444_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0218_),
    .Q(\as1802.regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7445_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0219_),
    .Q(\as1802.regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7446_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net670),
    .Q(\as1802.regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7447_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0221_),
    .Q(\as1802.regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7448_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0222_),
    .Q(\as1802.regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7449_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net636),
    .Q(\as1802.regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7450_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0224_),
    .Q(\as1802.regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7451_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0225_),
    .Q(\as1802.regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_4 _7452_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net285),
    .Q(_0008_));
 sky130_fd_sc_hd__dfxtp_4 _7453_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net743),
    .Q(_0009_));
 sky130_fd_sc_hd__dfxtp_2 _7454_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net777),
    .Q(_0010_));
 sky130_fd_sc_hd__dfxtp_2 _7455_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net311),
    .Q(_0011_));
 sky130_fd_sc_hd__dfxtp_1 _7456_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0226_),
    .Q(\as1802.regs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7457_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0227_),
    .Q(\as1802.regs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7458_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0228_),
    .Q(\as1802.regs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7459_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0229_),
    .Q(\as1802.regs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7460_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0230_),
    .Q(\as1802.regs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7461_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0231_),
    .Q(\as1802.regs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7462_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0232_),
    .Q(\as1802.regs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7463_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0233_),
    .Q(\as1802.regs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7464_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0234_),
    .Q(\as1802.regs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7465_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0235_),
    .Q(\as1802.regs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7466_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0236_),
    .Q(\as1802.regs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7467_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0237_),
    .Q(\as1802.regs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7468_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0238_),
    .Q(\as1802.regs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7469_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0239_),
    .Q(\as1802.regs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7470_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0240_),
    .Q(\as1802.regs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7471_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0241_),
    .Q(\as1802.regs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7472_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net734),
    .Q(\as1802.instr_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7473_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0013_),
    .Q(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7474_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_0014_),
    .Q(\as1802.instr_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7475_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net275),
    .Q(\as1802.instr_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7476_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0242_),
    .Q(\as1802.regs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7477_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0243_),
    .Q(\as1802.regs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7478_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0244_),
    .Q(\as1802.regs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7479_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0245_),
    .Q(\as1802.regs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7480_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0246_),
    .Q(\as1802.regs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7481_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0247_),
    .Q(\as1802.regs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7482_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0248_),
    .Q(\as1802.regs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7483_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0249_),
    .Q(\as1802.regs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7484_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0250_),
    .Q(\as1802.regs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7485_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0251_),
    .Q(\as1802.regs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7486_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0252_),
    .Q(\as1802.regs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7487_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0253_),
    .Q(\as1802.regs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7488_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0254_),
    .Q(\as1802.regs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7489_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0255_),
    .Q(\as1802.regs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7490_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0256_),
    .Q(\as1802.regs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7491_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0257_),
    .Q(\as1802.regs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7492_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net295),
    .Q(\as1802.MHI[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7493_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net301),
    .Q(\as1802.MHI[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7494_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net727),
    .Q(\as1802.MHI[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7495_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net305),
    .Q(\as1802.MHI[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7496_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net309),
    .Q(\as1802.MHI[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7497_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net320),
    .Q(\as1802.MHI[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7498_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net297),
    .Q(\as1802.MHI[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7499_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net376),
    .Q(\as1802.MHI[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7500_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net368),
    .Q(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7501_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net353),
    .Q(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7502_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0268_),
    .Q(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7503_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(net273),
    .Q(\as1802.addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7504_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net269),
    .Q(\as1802.addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7505_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net267),
    .Q(\as1802.addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7506_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net265),
    .Q(\as1802.addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7507_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net263),
    .Q(\as1802.addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7508_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(net257),
    .Q(\as1802.addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7509_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net259),
    .Q(\as1802.addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7510_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net261),
    .Q(\as1802.addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7511_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net293),
    .Q(\as1802.addr_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7512_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net291),
    .Q(\as1802.addr_buff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7513_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net303),
    .Q(\as1802.addr_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7514_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net283),
    .Q(\as1802.addr_buff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7515_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net299),
    .Q(\as1802.addr_buff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7516_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net287),
    .Q(\as1802.addr_buff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7517_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net281),
    .Q(\as1802.addr_buff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7518_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net307),
    .Q(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__dfxtp_2 _7519_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net399),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_2 _7520_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net393),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _7521_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net380),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _7522_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net365),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _7523_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net719),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_2 _7524_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net337),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_2 _7525_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net363),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _7526_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net386),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _7527_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net811),
    .Q(\as1802.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7528_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net330),
    .Q(\as1802.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7529_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0295_),
    .Q(\as1802.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7530_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net473),
    .Q(\as1802.X[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7531_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0297_),
    .Q(\as1802.last_hi_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7532_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0298_),
    .Q(\as1802.last_hi_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7533_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0299_),
    .Q(\as1802.last_hi_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7534_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0300_),
    .Q(\as1802.last_hi_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7535_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0301_),
    .Q(\as1802.last_hi_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7536_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_0302_),
    .Q(\as1802.last_hi_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7537_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0303_),
    .Q(\as1802.last_hi_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7538_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0304_),
    .Q(\as1802.last_hi_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7539_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(net832),
    .Q(\as1802.will_interrupt ));
 sky130_fd_sc_hd__dfxtp_4 _7540_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_0306_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _7541_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(net271),
    .Q(\as1802.MRD ));
 sky130_fd_sc_hd__dfxtp_4 _7542_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_0308_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_4 _7543_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(net339),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _7544_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0024_),
    .Q(\as1802.EF_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7545_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0025_),
    .Q(\as1802.EF_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7546_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0026_),
    .Q(\as1802.EF_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7547_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0027_),
    .Q(\as1802.EF_l[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7548_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0310_),
    .Q(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7549_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0311_),
    .Q(\as1802.instr_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7550_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0312_),
    .Q(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7551_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0313_),
    .Q(\as1802.cond_inv ));
 sky130_fd_sc_hd__dfxtp_1 _7552_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0314_),
    .Q(\as1802.instr_latch[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7553_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0315_),
    .Q(\as1802.instr_latch[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7554_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0316_),
    .Q(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7555_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0317_),
    .Q(\as1802.instr_latch[7] ));
 sky130_fd_sc_hd__dfxtp_4 _7556_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0318_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_4 _7557_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0319_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_4 _7558_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_0320_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_4 _7559_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(net835),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _7560_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0322_),
    .Q(\as1802.T[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7561_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0323_),
    .Q(\as1802.T[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7562_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0324_),
    .Q(\as1802.T[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7563_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0325_),
    .Q(\as1802.T[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7564_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0326_),
    .Q(\as1802.T[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7565_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0327_),
    .Q(\as1802.T[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7566_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0328_),
    .Q(\as1802.T[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7567_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0329_),
    .Q(\as1802.T[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7568_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net318),
    .Q(\as1802.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7569_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0331_),
    .Q(\as1802.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7570_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0332_),
    .Q(\as1802.P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7571_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0333_),
    .Q(\as1802.P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7572_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(net856),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _7573_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0335_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_2 _7574_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0336_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _7575_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(net850),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _7576_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(net877),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_2 _7577_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_0339_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _7578_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(net860),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _7579_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_0341_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_2 _7580_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net323),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_2 _7581_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net326),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_2 _7582_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net314),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _7583_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0345_),
    .Q(\as1802.D[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7584_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0346_),
    .Q(\as1802.D[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7585_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0347_),
    .Q(\as1802.D[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7586_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0348_),
    .Q(\as1802.D[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7587_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_0349_),
    .Q(\as1802.D[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7588_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0350_),
    .Q(\as1802.D[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7589_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0351_),
    .Q(\as1802.D[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7590_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_0352_),
    .Q(\as1802.D[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7591_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0353_),
    .Q(\as1802.regs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7592_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0354_),
    .Q(\as1802.regs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7593_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0355_),
    .Q(\as1802.regs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7594_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0356_),
    .Q(\as1802.regs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7595_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0357_),
    .Q(\as1802.regs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7596_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0358_),
    .Q(\as1802.regs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7597_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0359_),
    .Q(\as1802.regs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7598_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0360_),
    .Q(\as1802.regs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7599_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(net826),
    .Q(\as1802.mem_write ));
 sky130_fd_sc_hd__dfxtp_2 _7600_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0362_),
    .Q(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _7601_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0363_),
    .Q(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7602_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0364_),
    .Q(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7603_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net846),
    .Q(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _7604_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0366_),
    .Q(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7605_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0367_),
    .Q(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7606_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net870),
    .Q(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _7607_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net864),
    .Q(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7608_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0370_),
    .Q(\as1802.regs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7609_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0371_),
    .Q(\as1802.regs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7610_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0372_),
    .Q(\as1802.regs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7611_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0373_),
    .Q(\as1802.regs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7612_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0374_),
    .Q(\as1802.regs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7613_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0375_),
    .Q(\as1802.regs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7614_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0376_),
    .Q(\as1802.regs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7615_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0377_),
    .Q(\as1802.regs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7616_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0378_),
    .Q(\as1802.regs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7617_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0379_),
    .Q(\as1802.regs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7618_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0380_),
    .Q(\as1802.regs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7619_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0381_),
    .Q(\as1802.regs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7620_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0382_),
    .Q(\as1802.regs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7621_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0383_),
    .Q(\as1802.regs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7622_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0384_),
    .Q(\as1802.regs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7623_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0385_),
    .Q(\as1802.regs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7624_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net277),
    .Q(\as1802.lda ));
 sky130_fd_sc_hd__buf_1 _7630_ (.A(net21),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _7631_ (.A(net22),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_62_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(_0512_),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(_3503_),
    .X(net101));
 sky130_fd_sc_hd__buf_6 fanout102 (.A(_3483_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(_3483_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(_3482_),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(_3474_),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_3473_),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_8 fanout108 (.A(_3472_),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(_3472_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 fanout111 (.A(_3471_),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 fanout112 (.A(_3469_),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(_3469_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout114 (.A(_3467_),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout115 (.A(_3466_),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(_3466_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_8 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout118 (.A(_3443_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 fanout119 (.A(_3439_),
    .X(net119));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(net862),
    .X(net120));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(\as1802.D[7] ),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net861),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net853),
    .X(net126));
 sky130_fd_sc_hd__buf_6 fanout127 (.A(net881),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(\as1802.D[4] ),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(net872),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net875),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(net858),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(\as1802.D[1] ),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(net880),
    .X(net135));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(\as1802.D[0] ),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_6 fanout139 (.A(net55),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net142),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_8 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net54),
    .X(net142));
 sky130_fd_sc_hd__buf_8 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_8 fanout145 (.A(net53),
    .X(net145));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(net52),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_6 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_8 fanout151 (.A(net51),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_8 fanout152 (.A(net50),
    .X(net152));
 sky130_fd_sc_hd__buf_6 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_8 fanout154 (.A(net50),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_6 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(net49),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_8 fanout158 (.A(net160),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_6 fanout160 (.A(net48),
    .X(net160));
 sky130_fd_sc_hd__buf_6 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net57),
    .X(net162));
 sky130_fd_sc_hd__buf_8 fanout163 (.A(net882),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(\as1802.cond_inv ),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(\as1802.cond_inv ),
    .X(net166));
 sky130_fd_sc_hd__buf_6 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net821),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(net327),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net732),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(net883),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(_0011_),
    .X(net175));
 sky130_fd_sc_hd__buf_6 fanout176 (.A(_0010_),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_6 fanout178 (.A(_0009_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_6 fanout180 (.A(_0009_),
    .X(net180));
 sky130_fd_sc_hd__buf_8 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_8 fanout182 (.A(_0008_),
    .X(net182));
 sky130_fd_sc_hd__buf_8 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(_0008_),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout185 (.A(_0002_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_6 fanout187 (.A(_0001_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(_0001_),
    .X(net189));
 sky130_fd_sc_hd__buf_8 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_8 fanout191 (.A(_0000_),
    .X(net191));
 sky130_fd_sc_hd__buf_8 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_8 fanout193 (.A(_0000_),
    .X(net193));
 sky130_fd_sc_hd__buf_6 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_8 fanout195 (.A(_0007_),
    .X(net195));
 sky130_fd_sc_hd__buf_8 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(_0006_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(_0005_),
    .X(net199));
 sky130_fd_sc_hd__buf_6 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_8 fanout201 (.A(_0005_),
    .X(net201));
 sky130_fd_sc_hd__buf_8 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(_0004_),
    .X(net203));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_8 fanout205 (.A(_0004_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(_3464_),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(net209),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_6 fanout211 (.A(net44),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net44),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net44),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout77 (.A(_2321_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 fanout78 (.A(_0677_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_8 fanout80 (.A(_0685_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_8 fanout81 (.A(_0684_),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(_0657_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_8 fanout83 (.A(_0627_),
    .X(net83));
 sky130_fd_sc_hd__buf_6 fanout84 (.A(_0688_),
    .X(net84));
 sky130_fd_sc_hd__buf_4 fanout85 (.A(_0688_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(_2326_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_8 fanout88 (.A(_2322_),
    .X(net88));
 sky130_fd_sc_hd__buf_4 fanout89 (.A(_0831_),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(_0831_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 fanout91 (.A(net93),
    .X(net91));
 sky130_fd_sc_hd__buf_4 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(_0583_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(_0527_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_8 fanout95 (.A(_3500_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_8 fanout96 (.A(_3527_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_8 fanout97 (.A(_3509_),
    .X(net97));
 sky130_fd_sc_hd__buf_2 fanout98 (.A(_3509_),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0330_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\as1802.MHI[5] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0263_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net64),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_2659_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0342_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net65),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_2661_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0343_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\as1802.instr_latch[1] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0600_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0601_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0294_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\as1802.last_hi_addr[6] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_2475_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\as1802.last_hi_addr[0] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_2469_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net75),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_2464_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0290_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net59),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0309_),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\as1802.last_hi_addr[5] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_2474_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\as1802.T[3] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_2616_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\as1802.T[4] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_2617_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\as1802.T[1] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_2614_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\as1802.T[7] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_2620_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\as1802.T[2] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_2615_),
    .X(net351));
 sky130_fd_sc_hd__buf_2 hold134 (.A(\as1802.mem_cycle[0] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0267_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\as1802.T[0] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_2613_),
    .X(net355));
 sky130_fd_sc_hd__buf_2 hold138 (.A(\as1802.mem_cycle[2] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_2479_),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\as1802.T[6] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_2619_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\as1802.T[5] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_2618_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net76),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0291_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net73),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0288_),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_4 hold148 (.A(\as1802.mem_write ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_2309_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0266_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\as1802.last_hi_addr[4] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_2473_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\as1802.last_hi_addr[1] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_2470_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\as1802.last_hi_addr[3] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_2472_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\as1802.MHI[7] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0265_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\as1802.last_hi_addr[7] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_2476_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net72),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0287_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\as1802.regs[5][5] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0115_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\as1802.regs[3][8] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_3416_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net47),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0292_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\as1802.regs[6][4] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_1444_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\as1802.regs[6][0] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_1348_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\as1802.regs[1][12] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net71),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0286_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\as1802.regs[3][7] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_1535_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\as1802.regs[3][13] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_3421_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net70),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0285_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\as1802.regs[6][11] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_1311_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\as1802.regs[5][6] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_1544_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\as1802.regs[8][7] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_1671_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\as1802.regs[1][14] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\as1802.regs[13][13] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_1699_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\as1802.regs[4][8] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_1584_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\as1802.regs[5][12] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\as1802.regs[5][11] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_1323_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\as1802.regs[9][6] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_1660_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\as1802.regs[5][7] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_1545_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\as1802.regs[1][9] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\as1802.regs[9][15] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\as1802.regs[10][6] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\as1802.regs[10][14] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\as1802.regs[1][8] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_3406_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\as1802.regs[13][11] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_1697_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\as1802.regs[9][0] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_1654_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\as1802.regs[1][4] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\as1802.regs[6][12] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\as1802.regs[5][14] ),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 hold213 (.A(\as1802.X[0] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0016_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\as1802.regs[10][15] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\as1802.regs[6][8] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_1308_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\as1802.regs[10][12] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\as1802.regs[1][10] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_3408_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\as1802.regs[5][9] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\as1802.regs[4][11] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_1587_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\as1802.regs[6][9] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\as1802.regs[8][10] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_1288_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\as1802.regs[3][12] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\as1802.regs[0][9] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\as1802.regs[4][14] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\as1802.regs[9][11] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_3383_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\as1802.regs[8][6] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_1670_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\as1802.regs[10][0] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_1634_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\as1802.regs[1][11] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_3409_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\as1802.regs[8][2] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_1666_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0212_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\as1802.regs[6][14] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\as1802.regs[9][14] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\as1802.last_hi_addr[2] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_2471_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\as1802.regs[9][12] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\as1802.regs[6][13] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_1313_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\as1802.regs[12][8] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_1704_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\as1802.regs[4][5] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0099_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\as1802.regs[3][4] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_1532_),
    .X(net471));
 sky130_fd_sc_hd__buf_1 hold254 (.A(\as1802.X[3] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0296_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\as1802.regs[4][3] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\as1802.regs[13][2] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_1606_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0164_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\as1802.regs[4][6] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_1524_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\as1802.regs[8][11] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_1289_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\as1802.regs[10][8] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_1262_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\as1802.regs[3][15] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\as1802.regs[11][15] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\as1802.regs[9][2] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_1656_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0204_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\as1802.regs[4][9] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\as1802.regs[5][10] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_1322_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\as1802.regs[11][2] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_1626_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0180_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\as1802.regs[1][1] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_1559_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\as1802.regs[3][6] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\as1802.regs[6][10] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_1310_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\as1802.regs[7][4] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_1678_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\as1802.regs[9][5] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0207_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\as1802.regs[10][1] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_1635_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\as1802.regs[10][7] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_1641_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\as1802.regs[3][10] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_3418_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\as1802.regs[15][7] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_1601_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\as1802.regs[9][1] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_1655_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\as1802.regs[12][11] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_1707_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\as1802.regs[5][3] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\as1802.regs[4][7] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_1525_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\as1802.regs[13][15] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\as1802.regs[11][12] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\as1802.regs[9][7] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_1661_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\as1802.regs[13][14] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\as1802.regs[1][15] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\as1802.regs[0][10] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_1278_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\as1802.regs[4][4] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_1522_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\as1802.regs[9][10] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_3382_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\as1802.regs[8][13] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_1291_),
    .X(net532));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold315 (.A(net139),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0606_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0019_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\as1802.regs[10][4] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_1638_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\as1802.regs[4][0] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_1518_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\as1802.regs[4][15] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\as1802.regs[13][7] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_1611_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\as1802.regs[4][12] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\as1802.regs[15][6] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_1600_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\as1802.regs[7][9] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\as1802.regs[6][1] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_1370_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\as1802.regs[6][2] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\as1802.regs[5][4] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_1542_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\as1802.regs[10][2] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_1636_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0188_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\as1802.regs[8][3] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\as1802.regs[14][8] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_1684_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\as1802.regs[8][1] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_1665_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\as1802.regs[7][11] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_1301_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\as1802.regs[10][11] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_1265_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\as1802.regs[14][5] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0143_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\as1802.regs[0][13] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_1281_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\as1802.regs[1][13] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_3411_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\as1802.regs[0][8] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_1276_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\as1802.regs[7][0] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_1674_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\as1802.regs[15][2] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_1596_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0156_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\as1802.regs[5][0] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_1538_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\as1802.regs[13][4] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_1608_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\as1802.regs[0][14] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\as1802.regs[11][14] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\as1802.regs[1][6] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\as1802.regs[3][11] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_3419_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\as1802.regs[12][2] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_1616_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0172_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\as1802.regs[10][10] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_1264_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\as1802.regs[1][2] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\as1802.regs[12][7] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(_1621_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\as1802.regs[12][15] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\as1802.regs[3][1] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_1529_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\as1802.regs[8][15] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\as1802.addr_buff[5] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\as1802.regs[3][9] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\as1802.regs[12][5] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0175_),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\as1802.regs[12][6] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_1620_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\as1802.regs[8][9] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\as1802.regs[8][8] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_1286_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\as1802.regs[1][0] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_1558_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0274_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\as1802.regs[10][5] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0191_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\as1802.regs[7][13] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_1303_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\as1802.regs[0][1] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_1645_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\as1802.regs[12][14] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\as1802.regs[12][0] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_1614_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\as1802.regs[8][0] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\as1802.addr_buff[6] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_1664_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_0210_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\as1802.regs[13][3] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\as1802.regs[3][14] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\as1802.regs[0][5] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_0199_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\as1802.regs[7][14] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\as1802.regs[11][11] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_1717_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\as1802.regs[15][3] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0275_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\as1802.regs[14][10] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_1686_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\as1802.regs[3][2] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(_0104_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\as1802.regs[7][12] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\as1802.regs[13][5] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0167_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\as1802.regs[7][5] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0223_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\as1802.regs[8][5] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\as1802.addr_buff[7] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0215_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\as1802.regs[15][8] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0927_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\as1802.regs[6][6] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_1493_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\as1802.regs[7][8] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_1298_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\as1802.regs[12][12] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\as1802.regs[0][4] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_1648_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0276_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\as1802.regs[7][6] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_1680_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\as1802.regs[15][13] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_1166_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\as1802.regs[15][12] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\as1802.regs[11][13] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_1719_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\as1802.regs[13][10] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_1696_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\as1802.regs[11][10] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\as1802.addr_buff[4] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_1716_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\as1802.regs[11][9] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\as1802.regs[9][3] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\as1802.regs[15][4] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_1598_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\as1802.regs[0][12] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\as1802.regs[0][6] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\as1802.regs[15][11] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_1068_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\as1802.regs[12][10] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0273_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_1706_),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\as1802.regs[7][2] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0220_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\as1802.regs[12][9] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\as1802.regs[9][8] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_3380_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\as1802.regs[7][15] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\as1802.regs[10][9] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\as1802.regs[9][9] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\as1802.regs[12][13] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\as1802.addr_buff[3] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_1709_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\as1802.regs[14][15] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\as1802.regs[0][3] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\as1802.regs[14][9] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\as1802.regs[14][1] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_1575_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\as1802.regs[9][13] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_3385_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\as1802.regs[14][14] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\as1802.regs[0][11] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0272_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_1279_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\as1802.regs[15][14] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\as1802.regs[7][10] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_1300_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\as1802.regs[13][12] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\as1802.regs[8][14] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\as1802.regs[4][13] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_1589_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\as1802.regs[12][1] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_1615_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\as1802.addr_buff[2] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\as1802.regs[14][0] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_1574_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\as1802.regs[12][4] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_1618_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\as1802.regs[9][4] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_1658_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\as1802.regs[6][15] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\as1802.regs[0][0] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_1644_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\as1802.regs[4][10] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0271_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_1586_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\as1802.regs[0][7] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_1651_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\as1802.regs[5][13] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_1325_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\as1802.regs[0][15] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\as1802.regs[15][10] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_1023_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\as1802.regs[11][5] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(_0183_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\as1802.addr_buff[1] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net74),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0289_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\as1802.regs[14][2] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_1576_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0140_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\as1802.regs[11][6] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_1630_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0184_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\as1802.MHI[2] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_0260_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0270_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\as1802.regs[14][11] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_1687_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\as1802.regs[11][4] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_1628_),
    .X(net731));
 sky130_fd_sc_hd__buf_1 hold514 (.A(\as1802.instr_cycle[2] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0547_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0012_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\as1802.regs[12][3] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\as1802.regs[10][13] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_1267_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\as1802.MRD ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\as1802.regs[15][5] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0159_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\as1802.regs[10][3] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\as1802.regs[14][12] ),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_2 hold524 (.A(\as1802.P[1] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_0021_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\as1802.regs[13][0] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(_1604_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0162_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\as1802.regs[8][4] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0307_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_1668_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\as1802.regs[15][0] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_1594_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0154_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\as1802.regs[15][9] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\as1802.regs[11][7] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_1631_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\as1802.regs[13][1] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_1605_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\as1802.regs[11][1] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\as1802.addr_buff[0] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_1625_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\as1802.regs[1][5] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0131_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\as1802.regs[11][0] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_1624_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\as1802.regs[13][8] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_1694_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\as1802.regs[14][7] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_1581_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\as1802.regs[8][12] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0269_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\as1802.regs[4][2] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\as1802.regs[7][7] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_1681_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\as1802.regs[6][5] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0091_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\as1802.regs[3][0] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_1528_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\as1802.regs[5][2] ),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_2 hold558 (.A(\as1802.P[2] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0022_),
    .X(net777));
 sky130_fd_sc_hd__buf_1 hold56 (.A(\as1802.instr_cycle[3] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\as1802.regs[14][4] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_1578_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\as1802.regs[15][1] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_1595_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\as1802.regs[3][5] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_0107_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\as1802.regs[6][7] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(_1515_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\as1802.regs[1][7] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(_1565_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0015_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\as1802.regs[5][15] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\as1802.regs[13][9] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\as1802.regs[14][13] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_1689_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\as1802.regs[11][8] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(_1714_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\as1802.regs[6][3] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\as1802.regs[0][2] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\as1802.regs[5][8] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(_1320_),
    .X(net797));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold58 (.A(\as1802.lda ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\as1802.regs[5][1] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(_1539_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\as1802.regs[15][15] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\as1802.regs[1][3] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\as1802.regs[11][3] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\as1802.regs[14][6] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_1580_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(_0144_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\as1802.regs[13][6] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_1610_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0386_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0168_),
    .X(net808));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold591 (.A(\as1802.instr_latch[6] ),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_2 hold592 (.A(\as1802.instr_latch[0] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_0293_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\as1802.regs[7][1] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(_1675_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\as1802.regs[4][1] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(_1519_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\as1802.regs[14][3] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(net62),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_2 hold60 (.A(\as1802.X[1] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0037_),
    .X(net818));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold601 (.A(\as1802.X[2] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0018_),
    .X(net820));
 sky130_fd_sc_hd__buf_1 hold603 (.A(\as1802.instr_latch[2] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0605_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\as1802.regs[7][3] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\as1802.instr_cycle[1] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_3391_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0361_),
    .X(net826));
 sky130_fd_sc_hd__buf_1 hold609 (.A(\as1802.instr_latch[7] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0017_),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_2 hold610 (.A(net157),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\as1802.regs[3][3] ),
    .X(net829));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold612 (.A(\as1802.will_interrupt ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_2477_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0305_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(net46),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_2608_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_0321_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\as1802.regs[2][1] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_1549_),
    .X(net837));
 sky130_fd_sc_hd__buf_1 hold62 (.A(\as1802.addr_buff[14] ),
    .X(net280));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold620 (.A(\as1802.regs[2][13] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\as1802.regs[2][0] ),
    .X(net839));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold622 (.A(\as1802.regs[2][8] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\as1802.regs[2][6] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\as1802.regs[2][7] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\as1802.mem_cycle[1] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\as1802.regs[2][11] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_3399_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0365_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\as1802.regs[2][5] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0283_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0123_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(net151),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0337_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\as1802.regs[2][2] ),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 hold634 (.A(\as1802.instr_latch[5] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\as1802.D[5] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net60),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(net160),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0334_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\as1802.regs[2][3] ),
    .X(net857));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold64 (.A(\as1802.addr_buff[11] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\as1802.D[1] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(net142),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0340_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\as1802.D[6] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\as1802.D[7] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\as1802.regs[2][15] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0369_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(net67),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_2490_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\as1802.regs[2][9] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0280_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\as1802.regs[2][12] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\as1802.regs[2][14] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0368_),
    .X(net870));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold653 (.A(net63),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\as1802.D[3] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\as1802.regs[2][4] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\as1802.regs[2][10] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\as1802.D[2] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(net148),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_0338_),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_2 hold66 (.A(\as1802.P[0] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(net154),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net145),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\as1802.D[0] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\as1802.D[4] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\as1802.instr_latch[4] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\as1802.instr_cycle[0] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\as1802.regs[2][1] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(_1379_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\as1802.regs[2][13] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\as1802.instr_latch[2] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0020_),
    .X(net285));
 sky130_fd_sc_hd__buf_1 hold68 (.A(\as1802.addr_buff[13] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0282_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net61),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0036_),
    .X(net289));
 sky130_fd_sc_hd__buf_1 hold72 (.A(\as1802.addr_buff[9] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0278_),
    .X(net291));
 sky130_fd_sc_hd__buf_1 hold74 (.A(\as1802.addr_buff[8] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0277_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\as1802.MHI[0] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0258_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\as1802.MHI[6] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0264_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\as1802.P[3] ),
    .X(net890));
 sky130_fd_sc_hd__buf_1 hold80 (.A(\as1802.addr_buff[12] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0281_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\as1802.MHI[1] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0259_),
    .X(net301));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold84 (.A(\as1802.addr_buff[10] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0279_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\as1802.MHI[3] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0261_),
    .X(net305));
 sky130_fd_sc_hd__buf_1 hold88 (.A(\as1802.addr_buff[15] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0284_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\as1802.MHI[4] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0262_),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 hold92 (.A(net890),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0023_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net66),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_2663_),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0344_),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 hold97 (.A(\as1802.instr_latch[0] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0614_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0615_),
    .X(net317));
 sky130_fd_sc_hd__buf_1 input1 (.A(custom_settings[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(custom_settings[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(custom_settings[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(custom_settings[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(custom_settings[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(custom_settings[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(custom_settings[22]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(custom_settings[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(custom_settings[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(custom_settings[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(custom_settings[26]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(custom_settings[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(custom_settings[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(custom_settings[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(custom_settings[29]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(custom_settings[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(custom_settings[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(custom_settings[4]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(custom_settings[5]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(custom_settings[6]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(custom_settings[7]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(custom_settings[8]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(custom_settings[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(custom_settings[9]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(io_in[11]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(io_in[12]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(io_in[13]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(io_in[14]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(io_in[15]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(io_in[16]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(io_in[17]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(io_in[18]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(io_in[25]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(custom_settings[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(io_in[26]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(io_in[27]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(io_in[28]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(io_in[29]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(rst_n),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input5 (.A(custom_settings[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(custom_settings[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(custom_settings[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(custom_settings[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(custom_settings[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_oeb));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net159),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net156),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net154),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net150),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net148),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net242),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net141),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net138),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_1 output58 (.A(net58),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net61),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(io_out[35]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(io_out[9]));
 sky130_fd_sc_hd__buf_6 rebuffer1 (.A(_1764_),
    .X(net255));
 sky130_fd_sc_hd__buf_1 rebuffer10 (.A(_1938_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 rebuffer11 (.A(net228),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 rebuffer12 (.A(net234),
    .X(net230));
 sky130_fd_sc_hd__buf_6 rebuffer13 (.A(_3006_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 rebuffer14 (.A(net231),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 rebuffer16 (.A(_2834_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 rebuffer19 (.A(_1829_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 rebuffer2 (.A(_1900_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 rebuffer21 (.A(_1911_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(_1872_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(_1898_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(_1859_),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 rebuffer29 (.A(_1829_),
    .X(net247));
 sky130_fd_sc_hd__buf_1 rebuffer3 (.A(_1900_),
    .X(net221));
 sky130_fd_sc_hd__buf_6 rebuffer30 (.A(_1829_),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 rebuffer31 (.A(_1855_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 rebuffer33 (.A(_1829_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 rebuffer34 (.A(net888),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 rebuffer35 (.A(_1868_),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 rebuffer36 (.A(_1835_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_1856_),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(net252),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 rebuffer6 (.A(net223),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(_1916_),
    .X(net889));
 sky130_fd_sc_hd__buf_6 split1 (.A(_1829_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 split15 (.A(_2714_),
    .X(net233));
 sky130_fd_sc_hd__buf_1 split17 (.A(_3065_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 split18 (.A(_2874_),
    .X(net236));
 sky130_fd_sc_hd__buf_4 split20 (.A(net879),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 split24 (.A(net245),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 split25 (.A(_3012_),
    .X(net243));
 sky130_fd_sc_hd__buf_4 split26 (.A(net250),
    .X(net244));
 sky130_fd_sc_hd__dlymetal6s2s_1 split27 (.A(net144),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 split32 (.A(net143),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 split4 (.A(_3131_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 split7 (.A(_2948_),
    .X(net225));
 sky130_fd_sc_hd__buf_1 split8 (.A(_1722_),
    .X(net226));
 sky130_fd_sc_hd__buf_4 split9 (.A(_2838_),
    .X(net227));
 sky130_fd_sc_hd__buf_2 wire79 (.A(_2120_),
    .X(net79));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_218 (.LO(net218));
 assign io_out[25] = net214;
 assign io_out[26] = net215;
 assign io_out[27] = net216;
 assign io_out[28] = net217;
 assign io_out[29] = net218;
endmodule

