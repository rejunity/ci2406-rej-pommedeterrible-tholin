magic
tech sky130B
magscale 1 2
timestamp 1717499950
<< obsli1 >>
rect 1104 2159 38824 217617
<< obsm1 >>
rect 14 2128 39988 217648
<< metal2 >>
rect 2318 219200 2374 220000
rect 3054 219200 3110 220000
rect 3790 219200 3846 220000
rect 4526 219200 4582 220000
rect 5262 219200 5318 220000
rect 5998 219200 6054 220000
rect 6734 219200 6790 220000
rect 7470 219200 7526 220000
rect 8206 219200 8262 220000
rect 8942 219200 8998 220000
rect 9678 219200 9734 220000
rect 10414 219200 10470 220000
rect 11150 219200 11206 220000
rect 11886 219200 11942 220000
rect 12622 219200 12678 220000
rect 13358 219200 13414 220000
rect 14094 219200 14150 220000
rect 14830 219200 14886 220000
rect 15566 219200 15622 220000
rect 16302 219200 16358 220000
rect 17038 219200 17094 220000
rect 17774 219200 17830 220000
rect 18510 219200 18566 220000
rect 19246 219200 19302 220000
rect 19982 219200 20038 220000
rect 20718 219200 20774 220000
rect 21454 219200 21510 220000
rect 22190 219200 22246 220000
rect 22926 219200 22982 220000
rect 23662 219200 23718 220000
rect 24398 219200 24454 220000
rect 25134 219200 25190 220000
rect 25870 219200 25926 220000
rect 26606 219200 26662 220000
rect 27342 219200 27398 220000
rect 28078 219200 28134 220000
rect 28814 219200 28870 220000
rect 29550 219200 29606 220000
rect 30286 219200 30342 220000
rect 31022 219200 31078 220000
rect 31758 219200 31814 220000
rect 32494 219200 32550 220000
rect 33230 219200 33286 220000
rect 33966 219200 34022 220000
rect 34702 219200 34758 220000
rect 35438 219200 35494 220000
rect 36174 219200 36230 220000
rect 36910 219200 36966 220000
rect 37646 219200 37702 220000
rect 1122 0 1178 800
rect 2042 0 2098 800
rect 2962 0 3018 800
rect 3882 0 3938 800
rect 4802 0 4858 800
rect 5722 0 5778 800
rect 6642 0 6698 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 14002 0 14058 800
rect 14922 0 14978 800
rect 15842 0 15898 800
rect 16762 0 16818 800
rect 17682 0 17738 800
rect 18602 0 18658 800
rect 19522 0 19578 800
rect 20442 0 20498 800
rect 21362 0 21418 800
rect 22282 0 22338 800
rect 23202 0 23258 800
rect 24122 0 24178 800
rect 25042 0 25098 800
rect 25962 0 26018 800
rect 26882 0 26938 800
rect 27802 0 27858 800
rect 28722 0 28778 800
rect 29642 0 29698 800
rect 30562 0 30618 800
rect 31482 0 31538 800
rect 32402 0 32458 800
rect 33322 0 33378 800
rect 34242 0 34298 800
rect 35162 0 35218 800
rect 36082 0 36138 800
rect 37002 0 37058 800
rect 37922 0 37978 800
rect 38842 0 38898 800
<< obsm2 >>
rect 20 219144 2262 219314
rect 2430 219144 2998 219314
rect 3166 219144 3734 219314
rect 3902 219144 4470 219314
rect 4638 219144 5206 219314
rect 5374 219144 5942 219314
rect 6110 219144 6678 219314
rect 6846 219144 7414 219314
rect 7582 219144 8150 219314
rect 8318 219144 8886 219314
rect 9054 219144 9622 219314
rect 9790 219144 10358 219314
rect 10526 219144 11094 219314
rect 11262 219144 11830 219314
rect 11998 219144 12566 219314
rect 12734 219144 13302 219314
rect 13470 219144 14038 219314
rect 14206 219144 14774 219314
rect 14942 219144 15510 219314
rect 15678 219144 16246 219314
rect 16414 219144 16982 219314
rect 17150 219144 17718 219314
rect 17886 219144 18454 219314
rect 18622 219144 19190 219314
rect 19358 219144 19926 219314
rect 20094 219144 20662 219314
rect 20830 219144 21398 219314
rect 21566 219144 22134 219314
rect 22302 219144 22870 219314
rect 23038 219144 23606 219314
rect 23774 219144 24342 219314
rect 24510 219144 25078 219314
rect 25246 219144 25814 219314
rect 25982 219144 26550 219314
rect 26718 219144 27286 219314
rect 27454 219144 28022 219314
rect 28190 219144 28758 219314
rect 28926 219144 29494 219314
rect 29662 219144 30230 219314
rect 30398 219144 30966 219314
rect 31134 219144 31702 219314
rect 31870 219144 32438 219314
rect 32606 219144 33174 219314
rect 33342 219144 33910 219314
rect 34078 219144 34646 219314
rect 34814 219144 35382 219314
rect 35550 219144 36118 219314
rect 36286 219144 36854 219314
rect 37022 219144 37590 219314
rect 37758 219144 39988 219314
rect 20 856 39988 219144
rect 20 800 1066 856
rect 1234 800 1986 856
rect 2154 800 2906 856
rect 3074 800 3826 856
rect 3994 800 4746 856
rect 4914 800 5666 856
rect 5834 800 6586 856
rect 6754 800 7506 856
rect 7674 800 8426 856
rect 8594 800 9346 856
rect 9514 800 10266 856
rect 10434 800 11186 856
rect 11354 800 12106 856
rect 12274 800 13026 856
rect 13194 800 13946 856
rect 14114 800 14866 856
rect 15034 800 15786 856
rect 15954 800 16706 856
rect 16874 800 17626 856
rect 17794 800 18546 856
rect 18714 800 19466 856
rect 19634 800 20386 856
rect 20554 800 21306 856
rect 21474 800 22226 856
rect 22394 800 23146 856
rect 23314 800 24066 856
rect 24234 800 24986 856
rect 25154 800 25906 856
rect 26074 800 26826 856
rect 26994 800 27746 856
rect 27914 800 28666 856
rect 28834 800 29586 856
rect 29754 800 30506 856
rect 30674 800 31426 856
rect 31594 800 32346 856
rect 32514 800 33266 856
rect 33434 800 34186 856
rect 34354 800 35106 856
rect 35274 800 36026 856
rect 36194 800 36946 856
rect 37114 800 37866 856
rect 38034 800 38786 856
rect 38954 800 39988 856
<< metal3 >>
rect 0 199928 800 200048
rect 0 199112 800 199232
rect 0 198296 800 198416
rect 0 197480 800 197600
rect 0 196664 800 196784
rect 0 195848 800 195968
rect 0 195032 800 195152
rect 0 194216 800 194336
rect 0 193400 800 193520
rect 0 192584 800 192704
rect 0 191768 800 191888
rect 0 190952 800 191072
rect 0 190136 800 190256
rect 0 189320 800 189440
rect 39200 189320 40000 189440
rect 39200 188776 40000 188896
rect 0 188504 800 188624
rect 39200 188232 40000 188352
rect 0 187688 800 187808
rect 39200 187688 40000 187808
rect 39200 187144 40000 187264
rect 0 186872 800 186992
rect 39200 186600 40000 186720
rect 0 186056 800 186176
rect 39200 186056 40000 186176
rect 39200 185512 40000 185632
rect 0 185240 800 185360
rect 39200 184968 40000 185088
rect 0 184424 800 184544
rect 39200 184424 40000 184544
rect 39200 183880 40000 184000
rect 0 183608 800 183728
rect 39200 183336 40000 183456
rect 0 182792 800 182912
rect 39200 182792 40000 182912
rect 39200 182248 40000 182368
rect 0 181976 800 182096
rect 39200 181704 40000 181824
rect 0 181160 800 181280
rect 39200 181160 40000 181280
rect 39200 180616 40000 180736
rect 0 180344 800 180464
rect 39200 180072 40000 180192
rect 0 179528 800 179648
rect 39200 179528 40000 179648
rect 39200 178984 40000 179104
rect 0 178712 800 178832
rect 39200 178440 40000 178560
rect 0 177896 800 178016
rect 39200 177896 40000 178016
rect 39200 177352 40000 177472
rect 0 177080 800 177200
rect 39200 176808 40000 176928
rect 0 176264 800 176384
rect 39200 176264 40000 176384
rect 39200 175720 40000 175840
rect 0 175448 800 175568
rect 39200 175176 40000 175296
rect 0 174632 800 174752
rect 39200 174632 40000 174752
rect 39200 174088 40000 174208
rect 0 173816 800 173936
rect 39200 173544 40000 173664
rect 0 173000 800 173120
rect 39200 173000 40000 173120
rect 39200 172456 40000 172576
rect 0 172184 800 172304
rect 39200 171912 40000 172032
rect 0 171368 800 171488
rect 39200 171368 40000 171488
rect 39200 170824 40000 170944
rect 0 170552 800 170672
rect 39200 170280 40000 170400
rect 0 169736 800 169856
rect 39200 169736 40000 169856
rect 39200 169192 40000 169312
rect 0 168920 800 169040
rect 39200 168648 40000 168768
rect 0 168104 800 168224
rect 39200 168104 40000 168224
rect 39200 167560 40000 167680
rect 0 167288 800 167408
rect 39200 167016 40000 167136
rect 0 166472 800 166592
rect 39200 166472 40000 166592
rect 39200 165928 40000 166048
rect 0 165656 800 165776
rect 39200 165384 40000 165504
rect 0 164840 800 164960
rect 39200 164840 40000 164960
rect 39200 164296 40000 164416
rect 0 164024 800 164144
rect 39200 163752 40000 163872
rect 0 163208 800 163328
rect 39200 163208 40000 163328
rect 39200 162664 40000 162784
rect 0 162392 800 162512
rect 39200 162120 40000 162240
rect 0 161576 800 161696
rect 39200 161576 40000 161696
rect 39200 161032 40000 161152
rect 0 160760 800 160880
rect 39200 160488 40000 160608
rect 0 159944 800 160064
rect 39200 159944 40000 160064
rect 39200 159400 40000 159520
rect 0 159128 800 159248
rect 39200 158856 40000 158976
rect 0 158312 800 158432
rect 39200 158312 40000 158432
rect 39200 157768 40000 157888
rect 0 157496 800 157616
rect 39200 157224 40000 157344
rect 0 156680 800 156800
rect 39200 156680 40000 156800
rect 39200 156136 40000 156256
rect 0 155864 800 155984
rect 39200 155592 40000 155712
rect 0 155048 800 155168
rect 39200 155048 40000 155168
rect 39200 154504 40000 154624
rect 0 154232 800 154352
rect 39200 153960 40000 154080
rect 0 153416 800 153536
rect 39200 153416 40000 153536
rect 39200 152872 40000 152992
rect 0 152600 800 152720
rect 39200 152328 40000 152448
rect 0 151784 800 151904
rect 39200 151784 40000 151904
rect 39200 151240 40000 151360
rect 0 150968 800 151088
rect 39200 150696 40000 150816
rect 0 150152 800 150272
rect 39200 150152 40000 150272
rect 39200 149608 40000 149728
rect 0 149336 800 149456
rect 39200 149064 40000 149184
rect 0 148520 800 148640
rect 39200 148520 40000 148640
rect 39200 147976 40000 148096
rect 0 147704 800 147824
rect 39200 147432 40000 147552
rect 0 146888 800 147008
rect 39200 146888 40000 147008
rect 39200 146344 40000 146464
rect 0 146072 800 146192
rect 39200 145800 40000 145920
rect 0 145256 800 145376
rect 39200 145256 40000 145376
rect 39200 144712 40000 144832
rect 0 144440 800 144560
rect 39200 144168 40000 144288
rect 0 143624 800 143744
rect 39200 143624 40000 143744
rect 39200 143080 40000 143200
rect 0 142808 800 142928
rect 39200 142536 40000 142656
rect 0 141992 800 142112
rect 39200 141992 40000 142112
rect 39200 141448 40000 141568
rect 0 141176 800 141296
rect 39200 140904 40000 141024
rect 0 140360 800 140480
rect 39200 140360 40000 140480
rect 39200 139816 40000 139936
rect 0 139544 800 139664
rect 39200 139272 40000 139392
rect 0 138728 800 138848
rect 39200 138728 40000 138848
rect 39200 138184 40000 138304
rect 0 137912 800 138032
rect 39200 137640 40000 137760
rect 0 137096 800 137216
rect 39200 137096 40000 137216
rect 39200 136552 40000 136672
rect 0 136280 800 136400
rect 39200 136008 40000 136128
rect 0 135464 800 135584
rect 39200 135464 40000 135584
rect 39200 134920 40000 135040
rect 0 134648 800 134768
rect 39200 134376 40000 134496
rect 0 133832 800 133952
rect 39200 133832 40000 133952
rect 39200 133288 40000 133408
rect 0 133016 800 133136
rect 39200 132744 40000 132864
rect 0 132200 800 132320
rect 39200 132200 40000 132320
rect 39200 131656 40000 131776
rect 0 131384 800 131504
rect 39200 131112 40000 131232
rect 0 130568 800 130688
rect 39200 130568 40000 130688
rect 39200 130024 40000 130144
rect 0 129752 800 129872
rect 39200 129480 40000 129600
rect 0 128936 800 129056
rect 39200 128936 40000 129056
rect 39200 128392 40000 128512
rect 0 128120 800 128240
rect 39200 127848 40000 127968
rect 0 127304 800 127424
rect 39200 127304 40000 127424
rect 39200 126760 40000 126880
rect 0 126488 800 126608
rect 39200 126216 40000 126336
rect 0 125672 800 125792
rect 39200 125672 40000 125792
rect 39200 125128 40000 125248
rect 0 124856 800 124976
rect 39200 124584 40000 124704
rect 0 124040 800 124160
rect 39200 124040 40000 124160
rect 39200 123496 40000 123616
rect 0 123224 800 123344
rect 39200 122952 40000 123072
rect 0 122408 800 122528
rect 39200 122408 40000 122528
rect 39200 121864 40000 121984
rect 0 121592 800 121712
rect 39200 121320 40000 121440
rect 0 120776 800 120896
rect 39200 120776 40000 120896
rect 39200 120232 40000 120352
rect 0 119960 800 120080
rect 39200 119688 40000 119808
rect 0 119144 800 119264
rect 39200 119144 40000 119264
rect 39200 118600 40000 118720
rect 0 118328 800 118448
rect 39200 118056 40000 118176
rect 0 117512 800 117632
rect 39200 117512 40000 117632
rect 39200 116968 40000 117088
rect 0 116696 800 116816
rect 39200 116424 40000 116544
rect 0 115880 800 116000
rect 39200 115880 40000 116000
rect 39200 115336 40000 115456
rect 0 115064 800 115184
rect 39200 114792 40000 114912
rect 0 114248 800 114368
rect 39200 114248 40000 114368
rect 39200 113704 40000 113824
rect 0 113432 800 113552
rect 39200 113160 40000 113280
rect 0 112616 800 112736
rect 39200 112616 40000 112736
rect 39200 112072 40000 112192
rect 0 111800 800 111920
rect 39200 111528 40000 111648
rect 0 110984 800 111104
rect 39200 110984 40000 111104
rect 39200 110440 40000 110560
rect 0 110168 800 110288
rect 39200 109896 40000 110016
rect 0 109352 800 109472
rect 39200 109352 40000 109472
rect 39200 108808 40000 108928
rect 0 108536 800 108656
rect 39200 108264 40000 108384
rect 0 107720 800 107840
rect 39200 107720 40000 107840
rect 39200 107176 40000 107296
rect 0 106904 800 107024
rect 39200 106632 40000 106752
rect 0 106088 800 106208
rect 39200 106088 40000 106208
rect 39200 105544 40000 105664
rect 0 105272 800 105392
rect 39200 105000 40000 105120
rect 0 104456 800 104576
rect 39200 104456 40000 104576
rect 39200 103912 40000 104032
rect 0 103640 800 103760
rect 39200 103368 40000 103488
rect 0 102824 800 102944
rect 39200 102824 40000 102944
rect 39200 102280 40000 102400
rect 0 102008 800 102128
rect 39200 101736 40000 101856
rect 0 101192 800 101312
rect 39200 101192 40000 101312
rect 39200 100648 40000 100768
rect 0 100376 800 100496
rect 39200 100104 40000 100224
rect 0 99560 800 99680
rect 39200 99560 40000 99680
rect 39200 99016 40000 99136
rect 0 98744 800 98864
rect 39200 98472 40000 98592
rect 0 97928 800 98048
rect 39200 97928 40000 98048
rect 39200 97384 40000 97504
rect 0 97112 800 97232
rect 39200 96840 40000 96960
rect 0 96296 800 96416
rect 39200 96296 40000 96416
rect 39200 95752 40000 95872
rect 0 95480 800 95600
rect 39200 95208 40000 95328
rect 0 94664 800 94784
rect 39200 94664 40000 94784
rect 39200 94120 40000 94240
rect 0 93848 800 93968
rect 39200 93576 40000 93696
rect 0 93032 800 93152
rect 39200 93032 40000 93152
rect 39200 92488 40000 92608
rect 0 92216 800 92336
rect 39200 91944 40000 92064
rect 0 91400 800 91520
rect 39200 91400 40000 91520
rect 39200 90856 40000 90976
rect 0 90584 800 90704
rect 39200 90312 40000 90432
rect 0 89768 800 89888
rect 39200 89768 40000 89888
rect 39200 89224 40000 89344
rect 0 88952 800 89072
rect 39200 88680 40000 88800
rect 0 88136 800 88256
rect 39200 88136 40000 88256
rect 39200 87592 40000 87712
rect 0 87320 800 87440
rect 39200 87048 40000 87168
rect 0 86504 800 86624
rect 39200 86504 40000 86624
rect 39200 85960 40000 86080
rect 0 85688 800 85808
rect 39200 85416 40000 85536
rect 0 84872 800 84992
rect 39200 84872 40000 84992
rect 39200 84328 40000 84448
rect 0 84056 800 84176
rect 39200 83784 40000 83904
rect 0 83240 800 83360
rect 39200 83240 40000 83360
rect 39200 82696 40000 82816
rect 0 82424 800 82544
rect 39200 82152 40000 82272
rect 0 81608 800 81728
rect 39200 81608 40000 81728
rect 39200 81064 40000 81184
rect 0 80792 800 80912
rect 39200 80520 40000 80640
rect 0 79976 800 80096
rect 39200 79976 40000 80096
rect 39200 79432 40000 79552
rect 0 79160 800 79280
rect 39200 78888 40000 79008
rect 0 78344 800 78464
rect 39200 78344 40000 78464
rect 39200 77800 40000 77920
rect 0 77528 800 77648
rect 39200 77256 40000 77376
rect 0 76712 800 76832
rect 39200 76712 40000 76832
rect 39200 76168 40000 76288
rect 0 75896 800 76016
rect 39200 75624 40000 75744
rect 0 75080 800 75200
rect 39200 75080 40000 75200
rect 39200 74536 40000 74656
rect 0 74264 800 74384
rect 39200 73992 40000 74112
rect 0 73448 800 73568
rect 39200 73448 40000 73568
rect 39200 72904 40000 73024
rect 0 72632 800 72752
rect 39200 72360 40000 72480
rect 0 71816 800 71936
rect 39200 71816 40000 71936
rect 39200 71272 40000 71392
rect 0 71000 800 71120
rect 39200 70728 40000 70848
rect 0 70184 800 70304
rect 39200 70184 40000 70304
rect 39200 69640 40000 69760
rect 0 69368 800 69488
rect 39200 69096 40000 69216
rect 0 68552 800 68672
rect 39200 68552 40000 68672
rect 39200 68008 40000 68128
rect 0 67736 800 67856
rect 39200 67464 40000 67584
rect 0 66920 800 67040
rect 39200 66920 40000 67040
rect 39200 66376 40000 66496
rect 0 66104 800 66224
rect 39200 65832 40000 65952
rect 0 65288 800 65408
rect 39200 65288 40000 65408
rect 39200 64744 40000 64864
rect 0 64472 800 64592
rect 39200 64200 40000 64320
rect 0 63656 800 63776
rect 39200 63656 40000 63776
rect 39200 63112 40000 63232
rect 0 62840 800 62960
rect 39200 62568 40000 62688
rect 0 62024 800 62144
rect 39200 62024 40000 62144
rect 39200 61480 40000 61600
rect 0 61208 800 61328
rect 39200 60936 40000 61056
rect 0 60392 800 60512
rect 39200 60392 40000 60512
rect 39200 59848 40000 59968
rect 0 59576 800 59696
rect 39200 59304 40000 59424
rect 0 58760 800 58880
rect 39200 58760 40000 58880
rect 39200 58216 40000 58336
rect 0 57944 800 58064
rect 39200 57672 40000 57792
rect 0 57128 800 57248
rect 39200 57128 40000 57248
rect 39200 56584 40000 56704
rect 0 56312 800 56432
rect 39200 56040 40000 56160
rect 0 55496 800 55616
rect 39200 55496 40000 55616
rect 39200 54952 40000 55072
rect 0 54680 800 54800
rect 39200 54408 40000 54528
rect 0 53864 800 53984
rect 39200 53864 40000 53984
rect 39200 53320 40000 53440
rect 0 53048 800 53168
rect 39200 52776 40000 52896
rect 0 52232 800 52352
rect 39200 52232 40000 52352
rect 39200 51688 40000 51808
rect 0 51416 800 51536
rect 39200 51144 40000 51264
rect 0 50600 800 50720
rect 39200 50600 40000 50720
rect 39200 50056 40000 50176
rect 0 49784 800 49904
rect 39200 49512 40000 49632
rect 0 48968 800 49088
rect 39200 48968 40000 49088
rect 39200 48424 40000 48544
rect 0 48152 800 48272
rect 39200 47880 40000 48000
rect 0 47336 800 47456
rect 39200 47336 40000 47456
rect 39200 46792 40000 46912
rect 0 46520 800 46640
rect 39200 46248 40000 46368
rect 0 45704 800 45824
rect 39200 45704 40000 45824
rect 39200 45160 40000 45280
rect 0 44888 800 45008
rect 39200 44616 40000 44736
rect 0 44072 800 44192
rect 39200 44072 40000 44192
rect 39200 43528 40000 43648
rect 0 43256 800 43376
rect 39200 42984 40000 43104
rect 0 42440 800 42560
rect 39200 42440 40000 42560
rect 39200 41896 40000 42016
rect 0 41624 800 41744
rect 39200 41352 40000 41472
rect 0 40808 800 40928
rect 39200 40808 40000 40928
rect 39200 40264 40000 40384
rect 0 39992 800 40112
rect 39200 39720 40000 39840
rect 0 39176 800 39296
rect 39200 39176 40000 39296
rect 39200 38632 40000 38752
rect 0 38360 800 38480
rect 39200 38088 40000 38208
rect 0 37544 800 37664
rect 39200 37544 40000 37664
rect 39200 37000 40000 37120
rect 0 36728 800 36848
rect 39200 36456 40000 36576
rect 0 35912 800 36032
rect 39200 35912 40000 36032
rect 39200 35368 40000 35488
rect 0 35096 800 35216
rect 39200 34824 40000 34944
rect 0 34280 800 34400
rect 39200 34280 40000 34400
rect 39200 33736 40000 33856
rect 0 33464 800 33584
rect 39200 33192 40000 33312
rect 0 32648 800 32768
rect 39200 32648 40000 32768
rect 39200 32104 40000 32224
rect 0 31832 800 31952
rect 39200 31560 40000 31680
rect 0 31016 800 31136
rect 39200 31016 40000 31136
rect 39200 30472 40000 30592
rect 0 30200 800 30320
rect 0 29384 800 29504
rect 0 28568 800 28688
rect 0 27752 800 27872
rect 0 26936 800 27056
rect 0 26120 800 26240
rect 0 25304 800 25424
rect 0 24488 800 24608
rect 0 23672 800 23792
rect 0 22856 800 22976
rect 0 22040 800 22160
rect 0 21224 800 21344
rect 0 20408 800 20528
rect 0 19592 800 19712
<< obsm3 >>
rect 105 200128 39200 217633
rect 880 199848 39200 200128
rect 105 199312 39200 199848
rect 880 199032 39200 199312
rect 105 198496 39200 199032
rect 880 198216 39200 198496
rect 105 197680 39200 198216
rect 880 197400 39200 197680
rect 105 196864 39200 197400
rect 880 196584 39200 196864
rect 105 196048 39200 196584
rect 880 195768 39200 196048
rect 105 195232 39200 195768
rect 880 194952 39200 195232
rect 105 194416 39200 194952
rect 880 194136 39200 194416
rect 105 193600 39200 194136
rect 880 193320 39200 193600
rect 105 192784 39200 193320
rect 880 192504 39200 192784
rect 105 191968 39200 192504
rect 880 191688 39200 191968
rect 105 191152 39200 191688
rect 880 190872 39200 191152
rect 105 190336 39200 190872
rect 880 190056 39200 190336
rect 105 189520 39200 190056
rect 880 189240 39120 189520
rect 105 188976 39200 189240
rect 105 188704 39120 188976
rect 880 188696 39120 188704
rect 880 188432 39200 188696
rect 880 188424 39120 188432
rect 105 188152 39120 188424
rect 105 187888 39200 188152
rect 880 187608 39120 187888
rect 105 187344 39200 187608
rect 105 187072 39120 187344
rect 880 187064 39120 187072
rect 880 186800 39200 187064
rect 880 186792 39120 186800
rect 105 186520 39120 186792
rect 105 186256 39200 186520
rect 880 185976 39120 186256
rect 105 185712 39200 185976
rect 105 185440 39120 185712
rect 880 185432 39120 185440
rect 880 185168 39200 185432
rect 880 185160 39120 185168
rect 105 184888 39120 185160
rect 105 184624 39200 184888
rect 880 184344 39120 184624
rect 105 184080 39200 184344
rect 105 183808 39120 184080
rect 880 183800 39120 183808
rect 880 183536 39200 183800
rect 880 183528 39120 183536
rect 105 183256 39120 183528
rect 105 182992 39200 183256
rect 880 182712 39120 182992
rect 105 182448 39200 182712
rect 105 182176 39120 182448
rect 880 182168 39120 182176
rect 880 181904 39200 182168
rect 880 181896 39120 181904
rect 105 181624 39120 181896
rect 105 181360 39200 181624
rect 880 181080 39120 181360
rect 105 180816 39200 181080
rect 105 180544 39120 180816
rect 880 180536 39120 180544
rect 880 180272 39200 180536
rect 880 180264 39120 180272
rect 105 179992 39120 180264
rect 105 179728 39200 179992
rect 880 179448 39120 179728
rect 105 179184 39200 179448
rect 105 178912 39120 179184
rect 880 178904 39120 178912
rect 880 178640 39200 178904
rect 880 178632 39120 178640
rect 105 178360 39120 178632
rect 105 178096 39200 178360
rect 880 177816 39120 178096
rect 105 177552 39200 177816
rect 105 177280 39120 177552
rect 880 177272 39120 177280
rect 880 177008 39200 177272
rect 880 177000 39120 177008
rect 105 176728 39120 177000
rect 105 176464 39200 176728
rect 880 176184 39120 176464
rect 105 175920 39200 176184
rect 105 175648 39120 175920
rect 880 175640 39120 175648
rect 880 175376 39200 175640
rect 880 175368 39120 175376
rect 105 175096 39120 175368
rect 105 174832 39200 175096
rect 880 174552 39120 174832
rect 105 174288 39200 174552
rect 105 174016 39120 174288
rect 880 174008 39120 174016
rect 880 173744 39200 174008
rect 880 173736 39120 173744
rect 105 173464 39120 173736
rect 105 173200 39200 173464
rect 880 172920 39120 173200
rect 105 172656 39200 172920
rect 105 172384 39120 172656
rect 880 172376 39120 172384
rect 880 172112 39200 172376
rect 880 172104 39120 172112
rect 105 171832 39120 172104
rect 105 171568 39200 171832
rect 880 171288 39120 171568
rect 105 171024 39200 171288
rect 105 170752 39120 171024
rect 880 170744 39120 170752
rect 880 170480 39200 170744
rect 880 170472 39120 170480
rect 105 170200 39120 170472
rect 105 169936 39200 170200
rect 880 169656 39120 169936
rect 105 169392 39200 169656
rect 105 169120 39120 169392
rect 880 169112 39120 169120
rect 880 168848 39200 169112
rect 880 168840 39120 168848
rect 105 168568 39120 168840
rect 105 168304 39200 168568
rect 880 168024 39120 168304
rect 105 167760 39200 168024
rect 105 167488 39120 167760
rect 880 167480 39120 167488
rect 880 167216 39200 167480
rect 880 167208 39120 167216
rect 105 166936 39120 167208
rect 105 166672 39200 166936
rect 880 166392 39120 166672
rect 105 166128 39200 166392
rect 105 165856 39120 166128
rect 880 165848 39120 165856
rect 880 165584 39200 165848
rect 880 165576 39120 165584
rect 105 165304 39120 165576
rect 105 165040 39200 165304
rect 880 164760 39120 165040
rect 105 164496 39200 164760
rect 105 164224 39120 164496
rect 880 164216 39120 164224
rect 880 163952 39200 164216
rect 880 163944 39120 163952
rect 105 163672 39120 163944
rect 105 163408 39200 163672
rect 880 163128 39120 163408
rect 105 162864 39200 163128
rect 105 162592 39120 162864
rect 880 162584 39120 162592
rect 880 162320 39200 162584
rect 880 162312 39120 162320
rect 105 162040 39120 162312
rect 105 161776 39200 162040
rect 880 161496 39120 161776
rect 105 161232 39200 161496
rect 105 160960 39120 161232
rect 880 160952 39120 160960
rect 880 160688 39200 160952
rect 880 160680 39120 160688
rect 105 160408 39120 160680
rect 105 160144 39200 160408
rect 880 159864 39120 160144
rect 105 159600 39200 159864
rect 105 159328 39120 159600
rect 880 159320 39120 159328
rect 880 159056 39200 159320
rect 880 159048 39120 159056
rect 105 158776 39120 159048
rect 105 158512 39200 158776
rect 880 158232 39120 158512
rect 105 157968 39200 158232
rect 105 157696 39120 157968
rect 880 157688 39120 157696
rect 880 157424 39200 157688
rect 880 157416 39120 157424
rect 105 157144 39120 157416
rect 105 156880 39200 157144
rect 880 156600 39120 156880
rect 105 156336 39200 156600
rect 105 156064 39120 156336
rect 880 156056 39120 156064
rect 880 155792 39200 156056
rect 880 155784 39120 155792
rect 105 155512 39120 155784
rect 105 155248 39200 155512
rect 880 154968 39120 155248
rect 105 154704 39200 154968
rect 105 154432 39120 154704
rect 880 154424 39120 154432
rect 880 154160 39200 154424
rect 880 154152 39120 154160
rect 105 153880 39120 154152
rect 105 153616 39200 153880
rect 880 153336 39120 153616
rect 105 153072 39200 153336
rect 105 152800 39120 153072
rect 880 152792 39120 152800
rect 880 152528 39200 152792
rect 880 152520 39120 152528
rect 105 152248 39120 152520
rect 105 151984 39200 152248
rect 880 151704 39120 151984
rect 105 151440 39200 151704
rect 105 151168 39120 151440
rect 880 151160 39120 151168
rect 880 150896 39200 151160
rect 880 150888 39120 150896
rect 105 150616 39120 150888
rect 105 150352 39200 150616
rect 880 150072 39120 150352
rect 105 149808 39200 150072
rect 105 149536 39120 149808
rect 880 149528 39120 149536
rect 880 149264 39200 149528
rect 880 149256 39120 149264
rect 105 148984 39120 149256
rect 105 148720 39200 148984
rect 880 148440 39120 148720
rect 105 148176 39200 148440
rect 105 147904 39120 148176
rect 880 147896 39120 147904
rect 880 147632 39200 147896
rect 880 147624 39120 147632
rect 105 147352 39120 147624
rect 105 147088 39200 147352
rect 880 146808 39120 147088
rect 105 146544 39200 146808
rect 105 146272 39120 146544
rect 880 146264 39120 146272
rect 880 146000 39200 146264
rect 880 145992 39120 146000
rect 105 145720 39120 145992
rect 105 145456 39200 145720
rect 880 145176 39120 145456
rect 105 144912 39200 145176
rect 105 144640 39120 144912
rect 880 144632 39120 144640
rect 880 144368 39200 144632
rect 880 144360 39120 144368
rect 105 144088 39120 144360
rect 105 143824 39200 144088
rect 880 143544 39120 143824
rect 105 143280 39200 143544
rect 105 143008 39120 143280
rect 880 143000 39120 143008
rect 880 142736 39200 143000
rect 880 142728 39120 142736
rect 105 142456 39120 142728
rect 105 142192 39200 142456
rect 880 141912 39120 142192
rect 105 141648 39200 141912
rect 105 141376 39120 141648
rect 880 141368 39120 141376
rect 880 141104 39200 141368
rect 880 141096 39120 141104
rect 105 140824 39120 141096
rect 105 140560 39200 140824
rect 880 140280 39120 140560
rect 105 140016 39200 140280
rect 105 139744 39120 140016
rect 880 139736 39120 139744
rect 880 139472 39200 139736
rect 880 139464 39120 139472
rect 105 139192 39120 139464
rect 105 138928 39200 139192
rect 880 138648 39120 138928
rect 105 138384 39200 138648
rect 105 138112 39120 138384
rect 880 138104 39120 138112
rect 880 137840 39200 138104
rect 880 137832 39120 137840
rect 105 137560 39120 137832
rect 105 137296 39200 137560
rect 880 137016 39120 137296
rect 105 136752 39200 137016
rect 105 136480 39120 136752
rect 880 136472 39120 136480
rect 880 136208 39200 136472
rect 880 136200 39120 136208
rect 105 135928 39120 136200
rect 105 135664 39200 135928
rect 880 135384 39120 135664
rect 105 135120 39200 135384
rect 105 134848 39120 135120
rect 880 134840 39120 134848
rect 880 134576 39200 134840
rect 880 134568 39120 134576
rect 105 134296 39120 134568
rect 105 134032 39200 134296
rect 880 133752 39120 134032
rect 105 133488 39200 133752
rect 105 133216 39120 133488
rect 880 133208 39120 133216
rect 880 132944 39200 133208
rect 880 132936 39120 132944
rect 105 132664 39120 132936
rect 105 132400 39200 132664
rect 880 132120 39120 132400
rect 105 131856 39200 132120
rect 105 131584 39120 131856
rect 880 131576 39120 131584
rect 880 131312 39200 131576
rect 880 131304 39120 131312
rect 105 131032 39120 131304
rect 105 130768 39200 131032
rect 880 130488 39120 130768
rect 105 130224 39200 130488
rect 105 129952 39120 130224
rect 880 129944 39120 129952
rect 880 129680 39200 129944
rect 880 129672 39120 129680
rect 105 129400 39120 129672
rect 105 129136 39200 129400
rect 880 128856 39120 129136
rect 105 128592 39200 128856
rect 105 128320 39120 128592
rect 880 128312 39120 128320
rect 880 128048 39200 128312
rect 880 128040 39120 128048
rect 105 127768 39120 128040
rect 105 127504 39200 127768
rect 880 127224 39120 127504
rect 105 126960 39200 127224
rect 105 126688 39120 126960
rect 880 126680 39120 126688
rect 880 126416 39200 126680
rect 880 126408 39120 126416
rect 105 126136 39120 126408
rect 105 125872 39200 126136
rect 880 125592 39120 125872
rect 105 125328 39200 125592
rect 105 125056 39120 125328
rect 880 125048 39120 125056
rect 880 124784 39200 125048
rect 880 124776 39120 124784
rect 105 124504 39120 124776
rect 105 124240 39200 124504
rect 880 123960 39120 124240
rect 105 123696 39200 123960
rect 105 123424 39120 123696
rect 880 123416 39120 123424
rect 880 123152 39200 123416
rect 880 123144 39120 123152
rect 105 122872 39120 123144
rect 105 122608 39200 122872
rect 880 122328 39120 122608
rect 105 122064 39200 122328
rect 105 121792 39120 122064
rect 880 121784 39120 121792
rect 880 121520 39200 121784
rect 880 121512 39120 121520
rect 105 121240 39120 121512
rect 105 120976 39200 121240
rect 880 120696 39120 120976
rect 105 120432 39200 120696
rect 105 120160 39120 120432
rect 880 120152 39120 120160
rect 880 119888 39200 120152
rect 880 119880 39120 119888
rect 105 119608 39120 119880
rect 105 119344 39200 119608
rect 880 119064 39120 119344
rect 105 118800 39200 119064
rect 105 118528 39120 118800
rect 880 118520 39120 118528
rect 880 118256 39200 118520
rect 880 118248 39120 118256
rect 105 117976 39120 118248
rect 105 117712 39200 117976
rect 880 117432 39120 117712
rect 105 117168 39200 117432
rect 105 116896 39120 117168
rect 880 116888 39120 116896
rect 880 116624 39200 116888
rect 880 116616 39120 116624
rect 105 116344 39120 116616
rect 105 116080 39200 116344
rect 880 115800 39120 116080
rect 105 115536 39200 115800
rect 105 115264 39120 115536
rect 880 115256 39120 115264
rect 880 114992 39200 115256
rect 880 114984 39120 114992
rect 105 114712 39120 114984
rect 105 114448 39200 114712
rect 880 114168 39120 114448
rect 105 113904 39200 114168
rect 105 113632 39120 113904
rect 880 113624 39120 113632
rect 880 113360 39200 113624
rect 880 113352 39120 113360
rect 105 113080 39120 113352
rect 105 112816 39200 113080
rect 880 112536 39120 112816
rect 105 112272 39200 112536
rect 105 112000 39120 112272
rect 880 111992 39120 112000
rect 880 111728 39200 111992
rect 880 111720 39120 111728
rect 105 111448 39120 111720
rect 105 111184 39200 111448
rect 880 110904 39120 111184
rect 105 110640 39200 110904
rect 105 110368 39120 110640
rect 880 110360 39120 110368
rect 880 110096 39200 110360
rect 880 110088 39120 110096
rect 105 109816 39120 110088
rect 105 109552 39200 109816
rect 880 109272 39120 109552
rect 105 109008 39200 109272
rect 105 108736 39120 109008
rect 880 108728 39120 108736
rect 880 108464 39200 108728
rect 880 108456 39120 108464
rect 105 108184 39120 108456
rect 105 107920 39200 108184
rect 880 107640 39120 107920
rect 105 107376 39200 107640
rect 105 107104 39120 107376
rect 880 107096 39120 107104
rect 880 106832 39200 107096
rect 880 106824 39120 106832
rect 105 106552 39120 106824
rect 105 106288 39200 106552
rect 880 106008 39120 106288
rect 105 105744 39200 106008
rect 105 105472 39120 105744
rect 880 105464 39120 105472
rect 880 105200 39200 105464
rect 880 105192 39120 105200
rect 105 104920 39120 105192
rect 105 104656 39200 104920
rect 880 104376 39120 104656
rect 105 104112 39200 104376
rect 105 103840 39120 104112
rect 880 103832 39120 103840
rect 880 103568 39200 103832
rect 880 103560 39120 103568
rect 105 103288 39120 103560
rect 105 103024 39200 103288
rect 880 102744 39120 103024
rect 105 102480 39200 102744
rect 105 102208 39120 102480
rect 880 102200 39120 102208
rect 880 101936 39200 102200
rect 880 101928 39120 101936
rect 105 101656 39120 101928
rect 105 101392 39200 101656
rect 880 101112 39120 101392
rect 105 100848 39200 101112
rect 105 100576 39120 100848
rect 880 100568 39120 100576
rect 880 100304 39200 100568
rect 880 100296 39120 100304
rect 105 100024 39120 100296
rect 105 99760 39200 100024
rect 880 99480 39120 99760
rect 105 99216 39200 99480
rect 105 98944 39120 99216
rect 880 98936 39120 98944
rect 880 98672 39200 98936
rect 880 98664 39120 98672
rect 105 98392 39120 98664
rect 105 98128 39200 98392
rect 880 97848 39120 98128
rect 105 97584 39200 97848
rect 105 97312 39120 97584
rect 880 97304 39120 97312
rect 880 97040 39200 97304
rect 880 97032 39120 97040
rect 105 96760 39120 97032
rect 105 96496 39200 96760
rect 880 96216 39120 96496
rect 105 95952 39200 96216
rect 105 95680 39120 95952
rect 880 95672 39120 95680
rect 880 95408 39200 95672
rect 880 95400 39120 95408
rect 105 95128 39120 95400
rect 105 94864 39200 95128
rect 880 94584 39120 94864
rect 105 94320 39200 94584
rect 105 94048 39120 94320
rect 880 94040 39120 94048
rect 880 93776 39200 94040
rect 880 93768 39120 93776
rect 105 93496 39120 93768
rect 105 93232 39200 93496
rect 880 92952 39120 93232
rect 105 92688 39200 92952
rect 105 92416 39120 92688
rect 880 92408 39120 92416
rect 880 92144 39200 92408
rect 880 92136 39120 92144
rect 105 91864 39120 92136
rect 105 91600 39200 91864
rect 880 91320 39120 91600
rect 105 91056 39200 91320
rect 105 90784 39120 91056
rect 880 90776 39120 90784
rect 880 90512 39200 90776
rect 880 90504 39120 90512
rect 105 90232 39120 90504
rect 105 89968 39200 90232
rect 880 89688 39120 89968
rect 105 89424 39200 89688
rect 105 89152 39120 89424
rect 880 89144 39120 89152
rect 880 88880 39200 89144
rect 880 88872 39120 88880
rect 105 88600 39120 88872
rect 105 88336 39200 88600
rect 880 88056 39120 88336
rect 105 87792 39200 88056
rect 105 87520 39120 87792
rect 880 87512 39120 87520
rect 880 87248 39200 87512
rect 880 87240 39120 87248
rect 105 86968 39120 87240
rect 105 86704 39200 86968
rect 880 86424 39120 86704
rect 105 86160 39200 86424
rect 105 85888 39120 86160
rect 880 85880 39120 85888
rect 880 85616 39200 85880
rect 880 85608 39120 85616
rect 105 85336 39120 85608
rect 105 85072 39200 85336
rect 880 84792 39120 85072
rect 105 84528 39200 84792
rect 105 84256 39120 84528
rect 880 84248 39120 84256
rect 880 83984 39200 84248
rect 880 83976 39120 83984
rect 105 83704 39120 83976
rect 105 83440 39200 83704
rect 880 83160 39120 83440
rect 105 82896 39200 83160
rect 105 82624 39120 82896
rect 880 82616 39120 82624
rect 880 82352 39200 82616
rect 880 82344 39120 82352
rect 105 82072 39120 82344
rect 105 81808 39200 82072
rect 880 81528 39120 81808
rect 105 81264 39200 81528
rect 105 80992 39120 81264
rect 880 80984 39120 80992
rect 880 80720 39200 80984
rect 880 80712 39120 80720
rect 105 80440 39120 80712
rect 105 80176 39200 80440
rect 880 79896 39120 80176
rect 105 79632 39200 79896
rect 105 79360 39120 79632
rect 880 79352 39120 79360
rect 880 79088 39200 79352
rect 880 79080 39120 79088
rect 105 78808 39120 79080
rect 105 78544 39200 78808
rect 880 78264 39120 78544
rect 105 78000 39200 78264
rect 105 77728 39120 78000
rect 880 77720 39120 77728
rect 880 77456 39200 77720
rect 880 77448 39120 77456
rect 105 77176 39120 77448
rect 105 76912 39200 77176
rect 880 76632 39120 76912
rect 105 76368 39200 76632
rect 105 76096 39120 76368
rect 880 76088 39120 76096
rect 880 75824 39200 76088
rect 880 75816 39120 75824
rect 105 75544 39120 75816
rect 105 75280 39200 75544
rect 880 75000 39120 75280
rect 105 74736 39200 75000
rect 105 74464 39120 74736
rect 880 74456 39120 74464
rect 880 74192 39200 74456
rect 880 74184 39120 74192
rect 105 73912 39120 74184
rect 105 73648 39200 73912
rect 880 73368 39120 73648
rect 105 73104 39200 73368
rect 105 72832 39120 73104
rect 880 72824 39120 72832
rect 880 72560 39200 72824
rect 880 72552 39120 72560
rect 105 72280 39120 72552
rect 105 72016 39200 72280
rect 880 71736 39120 72016
rect 105 71472 39200 71736
rect 105 71200 39120 71472
rect 880 71192 39120 71200
rect 880 70928 39200 71192
rect 880 70920 39120 70928
rect 105 70648 39120 70920
rect 105 70384 39200 70648
rect 880 70104 39120 70384
rect 105 69840 39200 70104
rect 105 69568 39120 69840
rect 880 69560 39120 69568
rect 880 69296 39200 69560
rect 880 69288 39120 69296
rect 105 69016 39120 69288
rect 105 68752 39200 69016
rect 880 68472 39120 68752
rect 105 68208 39200 68472
rect 105 67936 39120 68208
rect 880 67928 39120 67936
rect 880 67664 39200 67928
rect 880 67656 39120 67664
rect 105 67384 39120 67656
rect 105 67120 39200 67384
rect 880 66840 39120 67120
rect 105 66576 39200 66840
rect 105 66304 39120 66576
rect 880 66296 39120 66304
rect 880 66032 39200 66296
rect 880 66024 39120 66032
rect 105 65752 39120 66024
rect 105 65488 39200 65752
rect 880 65208 39120 65488
rect 105 64944 39200 65208
rect 105 64672 39120 64944
rect 880 64664 39120 64672
rect 880 64400 39200 64664
rect 880 64392 39120 64400
rect 105 64120 39120 64392
rect 105 63856 39200 64120
rect 880 63576 39120 63856
rect 105 63312 39200 63576
rect 105 63040 39120 63312
rect 880 63032 39120 63040
rect 880 62768 39200 63032
rect 880 62760 39120 62768
rect 105 62488 39120 62760
rect 105 62224 39200 62488
rect 880 61944 39120 62224
rect 105 61680 39200 61944
rect 105 61408 39120 61680
rect 880 61400 39120 61408
rect 880 61136 39200 61400
rect 880 61128 39120 61136
rect 105 60856 39120 61128
rect 105 60592 39200 60856
rect 880 60312 39120 60592
rect 105 60048 39200 60312
rect 105 59776 39120 60048
rect 880 59768 39120 59776
rect 880 59504 39200 59768
rect 880 59496 39120 59504
rect 105 59224 39120 59496
rect 105 58960 39200 59224
rect 880 58680 39120 58960
rect 105 58416 39200 58680
rect 105 58144 39120 58416
rect 880 58136 39120 58144
rect 880 57872 39200 58136
rect 880 57864 39120 57872
rect 105 57592 39120 57864
rect 105 57328 39200 57592
rect 880 57048 39120 57328
rect 105 56784 39200 57048
rect 105 56512 39120 56784
rect 880 56504 39120 56512
rect 880 56240 39200 56504
rect 880 56232 39120 56240
rect 105 55960 39120 56232
rect 105 55696 39200 55960
rect 880 55416 39120 55696
rect 105 55152 39200 55416
rect 105 54880 39120 55152
rect 880 54872 39120 54880
rect 880 54608 39200 54872
rect 880 54600 39120 54608
rect 105 54328 39120 54600
rect 105 54064 39200 54328
rect 880 53784 39120 54064
rect 105 53520 39200 53784
rect 105 53248 39120 53520
rect 880 53240 39120 53248
rect 880 52976 39200 53240
rect 880 52968 39120 52976
rect 105 52696 39120 52968
rect 105 52432 39200 52696
rect 880 52152 39120 52432
rect 105 51888 39200 52152
rect 105 51616 39120 51888
rect 880 51608 39120 51616
rect 880 51344 39200 51608
rect 880 51336 39120 51344
rect 105 51064 39120 51336
rect 105 50800 39200 51064
rect 880 50520 39120 50800
rect 105 50256 39200 50520
rect 105 49984 39120 50256
rect 880 49976 39120 49984
rect 880 49712 39200 49976
rect 880 49704 39120 49712
rect 105 49432 39120 49704
rect 105 49168 39200 49432
rect 880 48888 39120 49168
rect 105 48624 39200 48888
rect 105 48352 39120 48624
rect 880 48344 39120 48352
rect 880 48080 39200 48344
rect 880 48072 39120 48080
rect 105 47800 39120 48072
rect 105 47536 39200 47800
rect 880 47256 39120 47536
rect 105 46992 39200 47256
rect 105 46720 39120 46992
rect 880 46712 39120 46720
rect 880 46448 39200 46712
rect 880 46440 39120 46448
rect 105 46168 39120 46440
rect 105 45904 39200 46168
rect 880 45624 39120 45904
rect 105 45360 39200 45624
rect 105 45088 39120 45360
rect 880 45080 39120 45088
rect 880 44816 39200 45080
rect 880 44808 39120 44816
rect 105 44536 39120 44808
rect 105 44272 39200 44536
rect 880 43992 39120 44272
rect 105 43728 39200 43992
rect 105 43456 39120 43728
rect 880 43448 39120 43456
rect 880 43184 39200 43448
rect 880 43176 39120 43184
rect 105 42904 39120 43176
rect 105 42640 39200 42904
rect 880 42360 39120 42640
rect 105 42096 39200 42360
rect 105 41824 39120 42096
rect 880 41816 39120 41824
rect 880 41552 39200 41816
rect 880 41544 39120 41552
rect 105 41272 39120 41544
rect 105 41008 39200 41272
rect 880 40728 39120 41008
rect 105 40464 39200 40728
rect 105 40192 39120 40464
rect 880 40184 39120 40192
rect 880 39920 39200 40184
rect 880 39912 39120 39920
rect 105 39640 39120 39912
rect 105 39376 39200 39640
rect 880 39096 39120 39376
rect 105 38832 39200 39096
rect 105 38560 39120 38832
rect 880 38552 39120 38560
rect 880 38288 39200 38552
rect 880 38280 39120 38288
rect 105 38008 39120 38280
rect 105 37744 39200 38008
rect 880 37464 39120 37744
rect 105 37200 39200 37464
rect 105 36928 39120 37200
rect 880 36920 39120 36928
rect 880 36656 39200 36920
rect 880 36648 39120 36656
rect 105 36376 39120 36648
rect 105 36112 39200 36376
rect 880 35832 39120 36112
rect 105 35568 39200 35832
rect 105 35296 39120 35568
rect 880 35288 39120 35296
rect 880 35024 39200 35288
rect 880 35016 39120 35024
rect 105 34744 39120 35016
rect 105 34480 39200 34744
rect 880 34200 39120 34480
rect 105 33936 39200 34200
rect 105 33664 39120 33936
rect 880 33656 39120 33664
rect 880 33392 39200 33656
rect 880 33384 39120 33392
rect 105 33112 39120 33384
rect 105 32848 39200 33112
rect 880 32568 39120 32848
rect 105 32304 39200 32568
rect 105 32032 39120 32304
rect 880 32024 39120 32032
rect 880 31760 39200 32024
rect 880 31752 39120 31760
rect 105 31480 39120 31752
rect 105 31216 39200 31480
rect 880 30936 39120 31216
rect 105 30672 39200 30936
rect 105 30400 39120 30672
rect 880 30392 39120 30400
rect 880 30120 39200 30392
rect 105 29584 39200 30120
rect 880 29304 39200 29584
rect 105 28768 39200 29304
rect 880 28488 39200 28768
rect 105 27952 39200 28488
rect 880 27672 39200 27952
rect 105 27136 39200 27672
rect 880 26856 39200 27136
rect 105 26320 39200 26856
rect 880 26040 39200 26320
rect 105 25504 39200 26040
rect 880 25224 39200 25504
rect 105 24688 39200 25224
rect 880 24408 39200 24688
rect 105 23872 39200 24408
rect 880 23592 39200 23872
rect 105 23056 39200 23592
rect 880 22776 39200 23056
rect 105 22240 39200 22776
rect 880 21960 39200 22240
rect 105 21424 39200 21960
rect 880 21144 39200 21424
rect 105 20608 39200 21144
rect 880 20328 39200 20608
rect 105 19792 39200 20328
rect 880 19512 39200 19792
rect 105 2143 39200 19512
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
<< obsm4 >>
rect 611 2755 4128 216069
rect 4608 2755 19488 216069
rect 19968 2755 34848 216069
rect 35328 2755 38213 216069
<< labels >>
rlabel metal2 s 31482 0 31538 800 6 cap_addr[0]
port 1 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 cap_addr[1]
port 2 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 cap_addr[2]
port 3 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 cap_addr[3]
port 4 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 cap_addr[4]
port 5 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 cap_addr[5]
port 6 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 cap_addr[6]
port 7 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 cap_addr[7]
port 8 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 cap_addr[8]
port 9 nsew signal output
rlabel metal2 s 3054 219200 3110 220000 6 cap_io_in[0]
port 10 nsew signal input
rlabel metal2 s 3790 219200 3846 220000 6 cap_io_in[1]
port 11 nsew signal input
rlabel metal2 s 4526 219200 4582 220000 6 cap_io_in[2]
port 12 nsew signal input
rlabel metal2 s 5262 219200 5318 220000 6 cap_io_in[3]
port 13 nsew signal input
rlabel metal2 s 5998 219200 6054 220000 6 cap_io_in[4]
port 14 nsew signal input
rlabel metal2 s 6734 219200 6790 220000 6 cap_io_in[5]
port 15 nsew signal input
rlabel metal2 s 7470 219200 7526 220000 6 cap_io_in[6]
port 16 nsew signal input
rlabel metal2 s 8206 219200 8262 220000 6 cap_io_in[7]
port 17 nsew signal input
rlabel metal2 s 8942 219200 8998 220000 6 cap_io_in[8]
port 18 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 custom_settings[0]
port 19 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 custom_settings[10]
port 20 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 custom_settings[11]
port 21 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 custom_settings[12]
port 22 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 custom_settings[13]
port 23 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 custom_settings[14]
port 24 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 custom_settings[15]
port 25 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 custom_settings[16]
port 26 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 custom_settings[17]
port 27 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 custom_settings[18]
port 28 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 custom_settings[19]
port 29 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 custom_settings[1]
port 30 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 custom_settings[20]
port 31 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 custom_settings[21]
port 32 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 custom_settings[22]
port 33 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 custom_settings[23]
port 34 nsew signal output
rlabel metal3 s 0 101192 800 101312 6 custom_settings[24]
port 35 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 custom_settings[25]
port 36 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 custom_settings[26]
port 37 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 custom_settings[27]
port 38 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 custom_settings[28]
port 39 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 custom_settings[29]
port 40 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 custom_settings[2]
port 41 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 custom_settings[30]
port 42 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 custom_settings[31]
port 43 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 custom_settings[3]
port 44 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 custom_settings[4]
port 45 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 custom_settings[5]
port 46 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 custom_settings[6]
port 47 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 custom_settings[7]
port 48 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 custom_settings[8]
port 49 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 custom_settings[9]
port 50 nsew signal output
rlabel metal2 s 2318 219200 2374 220000 6 io_in_0
port 51 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 io_oeb[0]
port 52 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 io_oeb[10]
port 53 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_oeb[11]
port 54 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 io_oeb[12]
port 55 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 io_oeb[13]
port 56 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 io_oeb[14]
port 57 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 io_oeb[15]
port 58 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 io_oeb[16]
port 59 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 io_oeb[17]
port 60 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 io_oeb[18]
port 61 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 io_oeb[19]
port 62 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 io_oeb[1]
port 63 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 io_oeb[20]
port 64 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_oeb[21]
port 65 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 io_oeb[22]
port 66 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 io_oeb[23]
port 67 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 io_oeb[24]
port 68 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 io_oeb[25]
port 69 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 io_oeb[26]
port 70 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 io_oeb[27]
port 71 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 io_oeb[28]
port 72 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 io_oeb[29]
port 73 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 io_oeb[2]
port 74 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 io_oeb[30]
port 75 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_oeb[31]
port 76 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 io_oeb[32]
port 77 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 io_oeb[33]
port 78 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 io_oeb[34]
port 79 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 io_oeb[35]
port 80 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 io_oeb[36]
port 81 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 io_oeb[37]
port 82 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_oeb[3]
port 83 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 io_oeb[4]
port 84 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 io_oeb[5]
port 85 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb[6]
port 86 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 io_oeb[7]
port 87 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[8]
port 88 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 io_oeb[9]
port 89 nsew signal output
rlabel metal3 s 39200 70728 40000 70848 6 io_oeb_6502
port 90 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 io_oeb_8x305[0]
port 91 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 io_oeb_8x305[1]
port 92 nsew signal input
rlabel metal3 s 0 197480 800 197600 6 io_oeb_8x305[2]
port 93 nsew signal input
rlabel metal3 s 0 198296 800 198416 6 io_oeb_8x305[3]
port 94 nsew signal input
rlabel metal3 s 0 199112 800 199232 6 io_oeb_8x305[4]
port 95 nsew signal input
rlabel metal3 s 39200 189320 40000 189440 6 io_oeb_as1802
port 96 nsew signal input
rlabel metal3 s 0 137096 800 137216 6 io_oeb_scrapcpu[0]
port 97 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 io_oeb_scrapcpu[10]
port 98 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 io_oeb_scrapcpu[11]
port 99 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 io_oeb_scrapcpu[12]
port 100 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 io_oeb_scrapcpu[13]
port 101 nsew signal input
rlabel metal3 s 0 148520 800 148640 6 io_oeb_scrapcpu[14]
port 102 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 io_oeb_scrapcpu[15]
port 103 nsew signal input
rlabel metal3 s 0 150152 800 150272 6 io_oeb_scrapcpu[16]
port 104 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 io_oeb_scrapcpu[17]
port 105 nsew signal input
rlabel metal3 s 0 151784 800 151904 6 io_oeb_scrapcpu[18]
port 106 nsew signal input
rlabel metal3 s 0 152600 800 152720 6 io_oeb_scrapcpu[19]
port 107 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 io_oeb_scrapcpu[1]
port 108 nsew signal input
rlabel metal3 s 0 153416 800 153536 6 io_oeb_scrapcpu[20]
port 109 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 io_oeb_scrapcpu[21]
port 110 nsew signal input
rlabel metal3 s 0 155048 800 155168 6 io_oeb_scrapcpu[22]
port 111 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 io_oeb_scrapcpu[23]
port 112 nsew signal input
rlabel metal3 s 0 156680 800 156800 6 io_oeb_scrapcpu[24]
port 113 nsew signal input
rlabel metal3 s 0 157496 800 157616 6 io_oeb_scrapcpu[25]
port 114 nsew signal input
rlabel metal3 s 0 158312 800 158432 6 io_oeb_scrapcpu[26]
port 115 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 io_oeb_scrapcpu[27]
port 116 nsew signal input
rlabel metal3 s 0 159944 800 160064 6 io_oeb_scrapcpu[28]
port 117 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 io_oeb_scrapcpu[29]
port 118 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 io_oeb_scrapcpu[2]
port 119 nsew signal input
rlabel metal3 s 0 161576 800 161696 6 io_oeb_scrapcpu[30]
port 120 nsew signal input
rlabel metal3 s 0 162392 800 162512 6 io_oeb_scrapcpu[31]
port 121 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 io_oeb_scrapcpu[32]
port 122 nsew signal input
rlabel metal3 s 0 164024 800 164144 6 io_oeb_scrapcpu[33]
port 123 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 io_oeb_scrapcpu[34]
port 124 nsew signal input
rlabel metal3 s 0 165656 800 165776 6 io_oeb_scrapcpu[35]
port 125 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 io_oeb_scrapcpu[3]
port 126 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 io_oeb_scrapcpu[4]
port 127 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 io_oeb_scrapcpu[5]
port 128 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 io_oeb_scrapcpu[6]
port 129 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 io_oeb_scrapcpu[7]
port 130 nsew signal input
rlabel metal3 s 0 143624 800 143744 6 io_oeb_scrapcpu[8]
port 131 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 io_oeb_scrapcpu[9]
port 132 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 io_oeb_vliw[0]
port 133 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 io_oeb_vliw[10]
port 134 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 io_oeb_vliw[11]
port 135 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 io_oeb_vliw[12]
port 136 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 io_oeb_vliw[13]
port 137 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 io_oeb_vliw[14]
port 138 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 io_oeb_vliw[15]
port 139 nsew signal input
rlabel metal3 s 0 120776 800 120896 6 io_oeb_vliw[16]
port 140 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 io_oeb_vliw[17]
port 141 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 io_oeb_vliw[18]
port 142 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 io_oeb_vliw[19]
port 143 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 io_oeb_vliw[1]
port 144 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 io_oeb_vliw[20]
port 145 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 io_oeb_vliw[21]
port 146 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 io_oeb_vliw[22]
port 147 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 io_oeb_vliw[23]
port 148 nsew signal input
rlabel metal3 s 0 127304 800 127424 6 io_oeb_vliw[24]
port 149 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 io_oeb_vliw[25]
port 150 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 io_oeb_vliw[26]
port 151 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 io_oeb_vliw[27]
port 152 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 io_oeb_vliw[28]
port 153 nsew signal input
rlabel metal3 s 0 131384 800 131504 6 io_oeb_vliw[29]
port 154 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 io_oeb_vliw[2]
port 155 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 io_oeb_vliw[30]
port 156 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 io_oeb_vliw[31]
port 157 nsew signal input
rlabel metal3 s 0 133832 800 133952 6 io_oeb_vliw[32]
port 158 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 io_oeb_vliw[33]
port 159 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 io_oeb_vliw[34]
port 160 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 io_oeb_vliw[35]
port 161 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 io_oeb_vliw[3]
port 162 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 io_oeb_vliw[4]
port 163 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 io_oeb_vliw[5]
port 164 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 io_oeb_vliw[6]
port 165 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 io_oeb_vliw[7]
port 166 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 io_oeb_vliw[8]
port 167 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 io_oeb_vliw[9]
port 168 nsew signal input
rlabel metal3 s 39200 130568 40000 130688 6 io_oeb_z80[0]
port 169 nsew signal input
rlabel metal3 s 39200 136008 40000 136128 6 io_oeb_z80[10]
port 170 nsew signal input
rlabel metal3 s 39200 136552 40000 136672 6 io_oeb_z80[11]
port 171 nsew signal input
rlabel metal3 s 39200 137096 40000 137216 6 io_oeb_z80[12]
port 172 nsew signal input
rlabel metal3 s 39200 137640 40000 137760 6 io_oeb_z80[13]
port 173 nsew signal input
rlabel metal3 s 39200 138184 40000 138304 6 io_oeb_z80[14]
port 174 nsew signal input
rlabel metal3 s 39200 138728 40000 138848 6 io_oeb_z80[15]
port 175 nsew signal input
rlabel metal3 s 39200 139272 40000 139392 6 io_oeb_z80[16]
port 176 nsew signal input
rlabel metal3 s 39200 139816 40000 139936 6 io_oeb_z80[17]
port 177 nsew signal input
rlabel metal3 s 39200 140360 40000 140480 6 io_oeb_z80[18]
port 178 nsew signal input
rlabel metal3 s 39200 140904 40000 141024 6 io_oeb_z80[19]
port 179 nsew signal input
rlabel metal3 s 39200 131112 40000 131232 6 io_oeb_z80[1]
port 180 nsew signal input
rlabel metal3 s 39200 141448 40000 141568 6 io_oeb_z80[20]
port 181 nsew signal input
rlabel metal3 s 39200 141992 40000 142112 6 io_oeb_z80[21]
port 182 nsew signal input
rlabel metal3 s 39200 142536 40000 142656 6 io_oeb_z80[22]
port 183 nsew signal input
rlabel metal3 s 39200 143080 40000 143200 6 io_oeb_z80[23]
port 184 nsew signal input
rlabel metal3 s 39200 143624 40000 143744 6 io_oeb_z80[24]
port 185 nsew signal input
rlabel metal3 s 39200 144168 40000 144288 6 io_oeb_z80[25]
port 186 nsew signal input
rlabel metal3 s 39200 144712 40000 144832 6 io_oeb_z80[26]
port 187 nsew signal input
rlabel metal3 s 39200 145256 40000 145376 6 io_oeb_z80[27]
port 188 nsew signal input
rlabel metal3 s 39200 145800 40000 145920 6 io_oeb_z80[28]
port 189 nsew signal input
rlabel metal3 s 39200 146344 40000 146464 6 io_oeb_z80[29]
port 190 nsew signal input
rlabel metal3 s 39200 131656 40000 131776 6 io_oeb_z80[2]
port 191 nsew signal input
rlabel metal3 s 39200 146888 40000 147008 6 io_oeb_z80[30]
port 192 nsew signal input
rlabel metal3 s 39200 147432 40000 147552 6 io_oeb_z80[31]
port 193 nsew signal input
rlabel metal3 s 39200 147976 40000 148096 6 io_oeb_z80[32]
port 194 nsew signal input
rlabel metal3 s 39200 148520 40000 148640 6 io_oeb_z80[33]
port 195 nsew signal input
rlabel metal3 s 39200 149064 40000 149184 6 io_oeb_z80[34]
port 196 nsew signal input
rlabel metal3 s 39200 149608 40000 149728 6 io_oeb_z80[35]
port 197 nsew signal input
rlabel metal3 s 39200 132200 40000 132320 6 io_oeb_z80[3]
port 198 nsew signal input
rlabel metal3 s 39200 132744 40000 132864 6 io_oeb_z80[4]
port 199 nsew signal input
rlabel metal3 s 39200 133288 40000 133408 6 io_oeb_z80[5]
port 200 nsew signal input
rlabel metal3 s 39200 133832 40000 133952 6 io_oeb_z80[6]
port 201 nsew signal input
rlabel metal3 s 39200 134376 40000 134496 6 io_oeb_z80[7]
port 202 nsew signal input
rlabel metal3 s 39200 134920 40000 135040 6 io_oeb_z80[8]
port 203 nsew signal input
rlabel metal3 s 39200 135464 40000 135584 6 io_oeb_z80[9]
port 204 nsew signal input
rlabel metal3 s 39200 30472 40000 30592 6 io_out[0]
port 205 nsew signal output
rlabel metal3 s 39200 35912 40000 36032 6 io_out[10]
port 206 nsew signal output
rlabel metal3 s 39200 36456 40000 36576 6 io_out[11]
port 207 nsew signal output
rlabel metal3 s 39200 37000 40000 37120 6 io_out[12]
port 208 nsew signal output
rlabel metal3 s 39200 37544 40000 37664 6 io_out[13]
port 209 nsew signal output
rlabel metal3 s 39200 38088 40000 38208 6 io_out[14]
port 210 nsew signal output
rlabel metal3 s 39200 38632 40000 38752 6 io_out[15]
port 211 nsew signal output
rlabel metal3 s 39200 39176 40000 39296 6 io_out[16]
port 212 nsew signal output
rlabel metal3 s 39200 39720 40000 39840 6 io_out[17]
port 213 nsew signal output
rlabel metal3 s 39200 40264 40000 40384 6 io_out[18]
port 214 nsew signal output
rlabel metal3 s 39200 40808 40000 40928 6 io_out[19]
port 215 nsew signal output
rlabel metal3 s 39200 31016 40000 31136 6 io_out[1]
port 216 nsew signal output
rlabel metal3 s 39200 41352 40000 41472 6 io_out[20]
port 217 nsew signal output
rlabel metal3 s 39200 41896 40000 42016 6 io_out[21]
port 218 nsew signal output
rlabel metal3 s 39200 42440 40000 42560 6 io_out[22]
port 219 nsew signal output
rlabel metal3 s 39200 42984 40000 43104 6 io_out[23]
port 220 nsew signal output
rlabel metal3 s 39200 43528 40000 43648 6 io_out[24]
port 221 nsew signal output
rlabel metal3 s 39200 44072 40000 44192 6 io_out[25]
port 222 nsew signal output
rlabel metal3 s 39200 44616 40000 44736 6 io_out[26]
port 223 nsew signal output
rlabel metal3 s 39200 45160 40000 45280 6 io_out[27]
port 224 nsew signal output
rlabel metal3 s 39200 45704 40000 45824 6 io_out[28]
port 225 nsew signal output
rlabel metal3 s 39200 46248 40000 46368 6 io_out[29]
port 226 nsew signal output
rlabel metal3 s 39200 31560 40000 31680 6 io_out[2]
port 227 nsew signal output
rlabel metal3 s 39200 46792 40000 46912 6 io_out[30]
port 228 nsew signal output
rlabel metal3 s 39200 47336 40000 47456 6 io_out[31]
port 229 nsew signal output
rlabel metal3 s 39200 47880 40000 48000 6 io_out[32]
port 230 nsew signal output
rlabel metal3 s 39200 48424 40000 48544 6 io_out[33]
port 231 nsew signal output
rlabel metal3 s 39200 48968 40000 49088 6 io_out[34]
port 232 nsew signal output
rlabel metal3 s 39200 49512 40000 49632 6 io_out[35]
port 233 nsew signal output
rlabel metal3 s 39200 50056 40000 50176 6 io_out[36]
port 234 nsew signal output
rlabel metal3 s 39200 50600 40000 50720 6 io_out[37]
port 235 nsew signal output
rlabel metal3 s 39200 32104 40000 32224 6 io_out[3]
port 236 nsew signal output
rlabel metal3 s 39200 32648 40000 32768 6 io_out[4]
port 237 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 io_out[5]
port 238 nsew signal output
rlabel metal3 s 39200 33736 40000 33856 6 io_out[6]
port 239 nsew signal output
rlabel metal3 s 39200 34280 40000 34400 6 io_out[7]
port 240 nsew signal output
rlabel metal3 s 39200 34824 40000 34944 6 io_out[8]
port 241 nsew signal output
rlabel metal3 s 39200 35368 40000 35488 6 io_out[9]
port 242 nsew signal output
rlabel metal3 s 39200 51144 40000 51264 6 io_out_6502[0]
port 243 nsew signal input
rlabel metal3 s 39200 56584 40000 56704 6 io_out_6502[10]
port 244 nsew signal input
rlabel metal3 s 39200 57128 40000 57248 6 io_out_6502[11]
port 245 nsew signal input
rlabel metal3 s 39200 57672 40000 57792 6 io_out_6502[12]
port 246 nsew signal input
rlabel metal3 s 39200 58216 40000 58336 6 io_out_6502[13]
port 247 nsew signal input
rlabel metal3 s 39200 58760 40000 58880 6 io_out_6502[14]
port 248 nsew signal input
rlabel metal3 s 39200 59304 40000 59424 6 io_out_6502[15]
port 249 nsew signal input
rlabel metal3 s 39200 59848 40000 59968 6 io_out_6502[16]
port 250 nsew signal input
rlabel metal3 s 39200 60392 40000 60512 6 io_out_6502[17]
port 251 nsew signal input
rlabel metal3 s 39200 60936 40000 61056 6 io_out_6502[18]
port 252 nsew signal input
rlabel metal3 s 39200 61480 40000 61600 6 io_out_6502[19]
port 253 nsew signal input
rlabel metal3 s 39200 51688 40000 51808 6 io_out_6502[1]
port 254 nsew signal input
rlabel metal3 s 39200 62024 40000 62144 6 io_out_6502[20]
port 255 nsew signal input
rlabel metal3 s 39200 62568 40000 62688 6 io_out_6502[21]
port 256 nsew signal input
rlabel metal3 s 39200 63112 40000 63232 6 io_out_6502[22]
port 257 nsew signal input
rlabel metal3 s 39200 63656 40000 63776 6 io_out_6502[23]
port 258 nsew signal input
rlabel metal3 s 39200 64200 40000 64320 6 io_out_6502[24]
port 259 nsew signal input
rlabel metal3 s 39200 64744 40000 64864 6 io_out_6502[25]
port 260 nsew signal input
rlabel metal3 s 39200 65288 40000 65408 6 io_out_6502[26]
port 261 nsew signal input
rlabel metal3 s 39200 65832 40000 65952 6 io_out_6502[27]
port 262 nsew signal input
rlabel metal3 s 39200 66376 40000 66496 6 io_out_6502[28]
port 263 nsew signal input
rlabel metal3 s 39200 66920 40000 67040 6 io_out_6502[29]
port 264 nsew signal input
rlabel metal3 s 39200 52232 40000 52352 6 io_out_6502[2]
port 265 nsew signal input
rlabel metal3 s 39200 67464 40000 67584 6 io_out_6502[30]
port 266 nsew signal input
rlabel metal3 s 39200 68008 40000 68128 6 io_out_6502[31]
port 267 nsew signal input
rlabel metal3 s 39200 68552 40000 68672 6 io_out_6502[32]
port 268 nsew signal input
rlabel metal3 s 39200 69096 40000 69216 6 io_out_6502[33]
port 269 nsew signal input
rlabel metal3 s 39200 69640 40000 69760 6 io_out_6502[34]
port 270 nsew signal input
rlabel metal3 s 39200 70184 40000 70304 6 io_out_6502[35]
port 271 nsew signal input
rlabel metal3 s 39200 52776 40000 52896 6 io_out_6502[3]
port 272 nsew signal input
rlabel metal3 s 39200 53320 40000 53440 6 io_out_6502[4]
port 273 nsew signal input
rlabel metal3 s 39200 53864 40000 53984 6 io_out_6502[5]
port 274 nsew signal input
rlabel metal3 s 39200 54408 40000 54528 6 io_out_6502[6]
port 275 nsew signal input
rlabel metal3 s 39200 54952 40000 55072 6 io_out_6502[7]
port 276 nsew signal input
rlabel metal3 s 39200 55496 40000 55616 6 io_out_6502[8]
port 277 nsew signal input
rlabel metal3 s 39200 56040 40000 56160 6 io_out_6502[9]
port 278 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 io_out_8x305[0]
port 279 nsew signal input
rlabel metal3 s 0 174632 800 174752 6 io_out_8x305[10]
port 280 nsew signal input
rlabel metal3 s 0 175448 800 175568 6 io_out_8x305[11]
port 281 nsew signal input
rlabel metal3 s 0 176264 800 176384 6 io_out_8x305[12]
port 282 nsew signal input
rlabel metal3 s 0 177080 800 177200 6 io_out_8x305[13]
port 283 nsew signal input
rlabel metal3 s 0 177896 800 178016 6 io_out_8x305[14]
port 284 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 io_out_8x305[15]
port 285 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 io_out_8x305[16]
port 286 nsew signal input
rlabel metal3 s 0 180344 800 180464 6 io_out_8x305[17]
port 287 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 io_out_8x305[18]
port 288 nsew signal input
rlabel metal3 s 0 181976 800 182096 6 io_out_8x305[19]
port 289 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 io_out_8x305[1]
port 290 nsew signal input
rlabel metal3 s 0 182792 800 182912 6 io_out_8x305[20]
port 291 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 io_out_8x305[21]
port 292 nsew signal input
rlabel metal3 s 0 184424 800 184544 6 io_out_8x305[22]
port 293 nsew signal input
rlabel metal3 s 0 185240 800 185360 6 io_out_8x305[23]
port 294 nsew signal input
rlabel metal3 s 0 186056 800 186176 6 io_out_8x305[24]
port 295 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 io_out_8x305[25]
port 296 nsew signal input
rlabel metal3 s 0 187688 800 187808 6 io_out_8x305[26]
port 297 nsew signal input
rlabel metal3 s 0 188504 800 188624 6 io_out_8x305[27]
port 298 nsew signal input
rlabel metal3 s 0 189320 800 189440 6 io_out_8x305[28]
port 299 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 io_out_8x305[29]
port 300 nsew signal input
rlabel metal3 s 0 168104 800 168224 6 io_out_8x305[2]
port 301 nsew signal input
rlabel metal3 s 0 190952 800 191072 6 io_out_8x305[30]
port 302 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 io_out_8x305[31]
port 303 nsew signal input
rlabel metal3 s 0 192584 800 192704 6 io_out_8x305[32]
port 304 nsew signal input
rlabel metal3 s 0 193400 800 193520 6 io_out_8x305[33]
port 305 nsew signal input
rlabel metal3 s 0 194216 800 194336 6 io_out_8x305[34]
port 306 nsew signal input
rlabel metal3 s 0 195032 800 195152 6 io_out_8x305[35]
port 307 nsew signal input
rlabel metal3 s 0 168920 800 169040 6 io_out_8x305[3]
port 308 nsew signal input
rlabel metal3 s 0 169736 800 169856 6 io_out_8x305[4]
port 309 nsew signal input
rlabel metal3 s 0 170552 800 170672 6 io_out_8x305[5]
port 310 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 io_out_8x305[6]
port 311 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 io_out_8x305[7]
port 312 nsew signal input
rlabel metal3 s 0 173000 800 173120 6 io_out_8x305[8]
port 313 nsew signal input
rlabel metal3 s 0 173816 800 173936 6 io_out_8x305[9]
port 314 nsew signal input
rlabel metal3 s 39200 169736 40000 169856 6 io_out_as1802[0]
port 315 nsew signal input
rlabel metal3 s 39200 175176 40000 175296 6 io_out_as1802[10]
port 316 nsew signal input
rlabel metal3 s 39200 175720 40000 175840 6 io_out_as1802[11]
port 317 nsew signal input
rlabel metal3 s 39200 176264 40000 176384 6 io_out_as1802[12]
port 318 nsew signal input
rlabel metal3 s 39200 176808 40000 176928 6 io_out_as1802[13]
port 319 nsew signal input
rlabel metal3 s 39200 177352 40000 177472 6 io_out_as1802[14]
port 320 nsew signal input
rlabel metal3 s 39200 177896 40000 178016 6 io_out_as1802[15]
port 321 nsew signal input
rlabel metal3 s 39200 178440 40000 178560 6 io_out_as1802[16]
port 322 nsew signal input
rlabel metal3 s 39200 178984 40000 179104 6 io_out_as1802[17]
port 323 nsew signal input
rlabel metal3 s 39200 179528 40000 179648 6 io_out_as1802[18]
port 324 nsew signal input
rlabel metal3 s 39200 180072 40000 180192 6 io_out_as1802[19]
port 325 nsew signal input
rlabel metal3 s 39200 170280 40000 170400 6 io_out_as1802[1]
port 326 nsew signal input
rlabel metal3 s 39200 180616 40000 180736 6 io_out_as1802[20]
port 327 nsew signal input
rlabel metal3 s 39200 181160 40000 181280 6 io_out_as1802[21]
port 328 nsew signal input
rlabel metal3 s 39200 181704 40000 181824 6 io_out_as1802[22]
port 329 nsew signal input
rlabel metal3 s 39200 182248 40000 182368 6 io_out_as1802[23]
port 330 nsew signal input
rlabel metal3 s 39200 182792 40000 182912 6 io_out_as1802[24]
port 331 nsew signal input
rlabel metal3 s 39200 183336 40000 183456 6 io_out_as1802[25]
port 332 nsew signal input
rlabel metal3 s 39200 183880 40000 184000 6 io_out_as1802[26]
port 333 nsew signal input
rlabel metal3 s 39200 184424 40000 184544 6 io_out_as1802[27]
port 334 nsew signal input
rlabel metal3 s 39200 184968 40000 185088 6 io_out_as1802[28]
port 335 nsew signal input
rlabel metal3 s 39200 185512 40000 185632 6 io_out_as1802[29]
port 336 nsew signal input
rlabel metal3 s 39200 170824 40000 170944 6 io_out_as1802[2]
port 337 nsew signal input
rlabel metal3 s 39200 186056 40000 186176 6 io_out_as1802[30]
port 338 nsew signal input
rlabel metal3 s 39200 186600 40000 186720 6 io_out_as1802[31]
port 339 nsew signal input
rlabel metal3 s 39200 187144 40000 187264 6 io_out_as1802[32]
port 340 nsew signal input
rlabel metal3 s 39200 187688 40000 187808 6 io_out_as1802[33]
port 341 nsew signal input
rlabel metal3 s 39200 188232 40000 188352 6 io_out_as1802[34]
port 342 nsew signal input
rlabel metal3 s 39200 188776 40000 188896 6 io_out_as1802[35]
port 343 nsew signal input
rlabel metal3 s 39200 171368 40000 171488 6 io_out_as1802[3]
port 344 nsew signal input
rlabel metal3 s 39200 171912 40000 172032 6 io_out_as1802[4]
port 345 nsew signal input
rlabel metal3 s 39200 172456 40000 172576 6 io_out_as1802[5]
port 346 nsew signal input
rlabel metal3 s 39200 173000 40000 173120 6 io_out_as1802[6]
port 347 nsew signal input
rlabel metal3 s 39200 173544 40000 173664 6 io_out_as1802[7]
port 348 nsew signal input
rlabel metal3 s 39200 174088 40000 174208 6 io_out_as1802[8]
port 349 nsew signal input
rlabel metal3 s 39200 174632 40000 174752 6 io_out_as1802[9]
port 350 nsew signal input
rlabel metal3 s 39200 150152 40000 150272 6 io_out_scrapcpu[0]
port 351 nsew signal input
rlabel metal3 s 39200 155592 40000 155712 6 io_out_scrapcpu[10]
port 352 nsew signal input
rlabel metal3 s 39200 156136 40000 156256 6 io_out_scrapcpu[11]
port 353 nsew signal input
rlabel metal3 s 39200 156680 40000 156800 6 io_out_scrapcpu[12]
port 354 nsew signal input
rlabel metal3 s 39200 157224 40000 157344 6 io_out_scrapcpu[13]
port 355 nsew signal input
rlabel metal3 s 39200 157768 40000 157888 6 io_out_scrapcpu[14]
port 356 nsew signal input
rlabel metal3 s 39200 158312 40000 158432 6 io_out_scrapcpu[15]
port 357 nsew signal input
rlabel metal3 s 39200 158856 40000 158976 6 io_out_scrapcpu[16]
port 358 nsew signal input
rlabel metal3 s 39200 159400 40000 159520 6 io_out_scrapcpu[17]
port 359 nsew signal input
rlabel metal3 s 39200 159944 40000 160064 6 io_out_scrapcpu[18]
port 360 nsew signal input
rlabel metal3 s 39200 160488 40000 160608 6 io_out_scrapcpu[19]
port 361 nsew signal input
rlabel metal3 s 39200 150696 40000 150816 6 io_out_scrapcpu[1]
port 362 nsew signal input
rlabel metal3 s 39200 161032 40000 161152 6 io_out_scrapcpu[20]
port 363 nsew signal input
rlabel metal3 s 39200 161576 40000 161696 6 io_out_scrapcpu[21]
port 364 nsew signal input
rlabel metal3 s 39200 162120 40000 162240 6 io_out_scrapcpu[22]
port 365 nsew signal input
rlabel metal3 s 39200 162664 40000 162784 6 io_out_scrapcpu[23]
port 366 nsew signal input
rlabel metal3 s 39200 163208 40000 163328 6 io_out_scrapcpu[24]
port 367 nsew signal input
rlabel metal3 s 39200 163752 40000 163872 6 io_out_scrapcpu[25]
port 368 nsew signal input
rlabel metal3 s 39200 164296 40000 164416 6 io_out_scrapcpu[26]
port 369 nsew signal input
rlabel metal3 s 39200 164840 40000 164960 6 io_out_scrapcpu[27]
port 370 nsew signal input
rlabel metal3 s 39200 165384 40000 165504 6 io_out_scrapcpu[28]
port 371 nsew signal input
rlabel metal3 s 39200 165928 40000 166048 6 io_out_scrapcpu[29]
port 372 nsew signal input
rlabel metal3 s 39200 151240 40000 151360 6 io_out_scrapcpu[2]
port 373 nsew signal input
rlabel metal3 s 39200 166472 40000 166592 6 io_out_scrapcpu[30]
port 374 nsew signal input
rlabel metal3 s 39200 167016 40000 167136 6 io_out_scrapcpu[31]
port 375 nsew signal input
rlabel metal3 s 39200 167560 40000 167680 6 io_out_scrapcpu[32]
port 376 nsew signal input
rlabel metal3 s 39200 168104 40000 168224 6 io_out_scrapcpu[33]
port 377 nsew signal input
rlabel metal3 s 39200 168648 40000 168768 6 io_out_scrapcpu[34]
port 378 nsew signal input
rlabel metal3 s 39200 169192 40000 169312 6 io_out_scrapcpu[35]
port 379 nsew signal input
rlabel metal3 s 39200 151784 40000 151904 6 io_out_scrapcpu[3]
port 380 nsew signal input
rlabel metal3 s 39200 152328 40000 152448 6 io_out_scrapcpu[4]
port 381 nsew signal input
rlabel metal3 s 39200 152872 40000 152992 6 io_out_scrapcpu[5]
port 382 nsew signal input
rlabel metal3 s 39200 153416 40000 153536 6 io_out_scrapcpu[6]
port 383 nsew signal input
rlabel metal3 s 39200 153960 40000 154080 6 io_out_scrapcpu[7]
port 384 nsew signal input
rlabel metal3 s 39200 154504 40000 154624 6 io_out_scrapcpu[8]
port 385 nsew signal input
rlabel metal3 s 39200 155048 40000 155168 6 io_out_scrapcpu[9]
port 386 nsew signal input
rlabel metal2 s 10414 219200 10470 220000 6 io_out_vliw[0]
port 387 nsew signal input
rlabel metal2 s 17774 219200 17830 220000 6 io_out_vliw[10]
port 388 nsew signal input
rlabel metal2 s 18510 219200 18566 220000 6 io_out_vliw[11]
port 389 nsew signal input
rlabel metal2 s 19246 219200 19302 220000 6 io_out_vliw[12]
port 390 nsew signal input
rlabel metal2 s 19982 219200 20038 220000 6 io_out_vliw[13]
port 391 nsew signal input
rlabel metal2 s 20718 219200 20774 220000 6 io_out_vliw[14]
port 392 nsew signal input
rlabel metal2 s 21454 219200 21510 220000 6 io_out_vliw[15]
port 393 nsew signal input
rlabel metal2 s 22190 219200 22246 220000 6 io_out_vliw[16]
port 394 nsew signal input
rlabel metal2 s 22926 219200 22982 220000 6 io_out_vliw[17]
port 395 nsew signal input
rlabel metal2 s 23662 219200 23718 220000 6 io_out_vliw[18]
port 396 nsew signal input
rlabel metal2 s 24398 219200 24454 220000 6 io_out_vliw[19]
port 397 nsew signal input
rlabel metal2 s 11150 219200 11206 220000 6 io_out_vliw[1]
port 398 nsew signal input
rlabel metal2 s 25134 219200 25190 220000 6 io_out_vliw[20]
port 399 nsew signal input
rlabel metal2 s 25870 219200 25926 220000 6 io_out_vliw[21]
port 400 nsew signal input
rlabel metal2 s 26606 219200 26662 220000 6 io_out_vliw[22]
port 401 nsew signal input
rlabel metal2 s 27342 219200 27398 220000 6 io_out_vliw[23]
port 402 nsew signal input
rlabel metal2 s 28078 219200 28134 220000 6 io_out_vliw[24]
port 403 nsew signal input
rlabel metal2 s 28814 219200 28870 220000 6 io_out_vliw[25]
port 404 nsew signal input
rlabel metal2 s 29550 219200 29606 220000 6 io_out_vliw[26]
port 405 nsew signal input
rlabel metal2 s 30286 219200 30342 220000 6 io_out_vliw[27]
port 406 nsew signal input
rlabel metal2 s 31022 219200 31078 220000 6 io_out_vliw[28]
port 407 nsew signal input
rlabel metal2 s 31758 219200 31814 220000 6 io_out_vliw[29]
port 408 nsew signal input
rlabel metal2 s 11886 219200 11942 220000 6 io_out_vliw[2]
port 409 nsew signal input
rlabel metal2 s 32494 219200 32550 220000 6 io_out_vliw[30]
port 410 nsew signal input
rlabel metal2 s 33230 219200 33286 220000 6 io_out_vliw[31]
port 411 nsew signal input
rlabel metal2 s 33966 219200 34022 220000 6 io_out_vliw[32]
port 412 nsew signal input
rlabel metal2 s 34702 219200 34758 220000 6 io_out_vliw[33]
port 413 nsew signal input
rlabel metal2 s 35438 219200 35494 220000 6 io_out_vliw[34]
port 414 nsew signal input
rlabel metal2 s 36174 219200 36230 220000 6 io_out_vliw[35]
port 415 nsew signal input
rlabel metal2 s 12622 219200 12678 220000 6 io_out_vliw[3]
port 416 nsew signal input
rlabel metal2 s 13358 219200 13414 220000 6 io_out_vliw[4]
port 417 nsew signal input
rlabel metal2 s 14094 219200 14150 220000 6 io_out_vliw[5]
port 418 nsew signal input
rlabel metal2 s 14830 219200 14886 220000 6 io_out_vliw[6]
port 419 nsew signal input
rlabel metal2 s 15566 219200 15622 220000 6 io_out_vliw[7]
port 420 nsew signal input
rlabel metal2 s 16302 219200 16358 220000 6 io_out_vliw[8]
port 421 nsew signal input
rlabel metal2 s 17038 219200 17094 220000 6 io_out_vliw[9]
port 422 nsew signal input
rlabel metal3 s 39200 110440 40000 110560 6 io_out_z80[0]
port 423 nsew signal input
rlabel metal3 s 39200 115880 40000 116000 6 io_out_z80[10]
port 424 nsew signal input
rlabel metal3 s 39200 116424 40000 116544 6 io_out_z80[11]
port 425 nsew signal input
rlabel metal3 s 39200 116968 40000 117088 6 io_out_z80[12]
port 426 nsew signal input
rlabel metal3 s 39200 117512 40000 117632 6 io_out_z80[13]
port 427 nsew signal input
rlabel metal3 s 39200 118056 40000 118176 6 io_out_z80[14]
port 428 nsew signal input
rlabel metal3 s 39200 118600 40000 118720 6 io_out_z80[15]
port 429 nsew signal input
rlabel metal3 s 39200 119144 40000 119264 6 io_out_z80[16]
port 430 nsew signal input
rlabel metal3 s 39200 119688 40000 119808 6 io_out_z80[17]
port 431 nsew signal input
rlabel metal3 s 39200 120232 40000 120352 6 io_out_z80[18]
port 432 nsew signal input
rlabel metal3 s 39200 120776 40000 120896 6 io_out_z80[19]
port 433 nsew signal input
rlabel metal3 s 39200 110984 40000 111104 6 io_out_z80[1]
port 434 nsew signal input
rlabel metal3 s 39200 121320 40000 121440 6 io_out_z80[20]
port 435 nsew signal input
rlabel metal3 s 39200 121864 40000 121984 6 io_out_z80[21]
port 436 nsew signal input
rlabel metal3 s 39200 122408 40000 122528 6 io_out_z80[22]
port 437 nsew signal input
rlabel metal3 s 39200 122952 40000 123072 6 io_out_z80[23]
port 438 nsew signal input
rlabel metal3 s 39200 123496 40000 123616 6 io_out_z80[24]
port 439 nsew signal input
rlabel metal3 s 39200 124040 40000 124160 6 io_out_z80[25]
port 440 nsew signal input
rlabel metal3 s 39200 124584 40000 124704 6 io_out_z80[26]
port 441 nsew signal input
rlabel metal3 s 39200 125128 40000 125248 6 io_out_z80[27]
port 442 nsew signal input
rlabel metal3 s 39200 125672 40000 125792 6 io_out_z80[28]
port 443 nsew signal input
rlabel metal3 s 39200 126216 40000 126336 6 io_out_z80[29]
port 444 nsew signal input
rlabel metal3 s 39200 111528 40000 111648 6 io_out_z80[2]
port 445 nsew signal input
rlabel metal3 s 39200 126760 40000 126880 6 io_out_z80[30]
port 446 nsew signal input
rlabel metal3 s 39200 127304 40000 127424 6 io_out_z80[31]
port 447 nsew signal input
rlabel metal3 s 39200 127848 40000 127968 6 io_out_z80[32]
port 448 nsew signal input
rlabel metal3 s 39200 128392 40000 128512 6 io_out_z80[33]
port 449 nsew signal input
rlabel metal3 s 39200 128936 40000 129056 6 io_out_z80[34]
port 450 nsew signal input
rlabel metal3 s 39200 129480 40000 129600 6 io_out_z80[35]
port 451 nsew signal input
rlabel metal3 s 39200 112072 40000 112192 6 io_out_z80[3]
port 452 nsew signal input
rlabel metal3 s 39200 112616 40000 112736 6 io_out_z80[4]
port 453 nsew signal input
rlabel metal3 s 39200 113160 40000 113280 6 io_out_z80[5]
port 454 nsew signal input
rlabel metal3 s 39200 113704 40000 113824 6 io_out_z80[6]
port 455 nsew signal input
rlabel metal3 s 39200 114248 40000 114368 6 io_out_z80[7]
port 456 nsew signal input
rlabel metal3 s 39200 114792 40000 114912 6 io_out_z80[8]
port 457 nsew signal input
rlabel metal3 s 39200 115336 40000 115456 6 io_out_z80[9]
port 458 nsew signal input
rlabel metal3 s 39200 88680 40000 88800 6 la_data_out[0]
port 459 nsew signal output
rlabel metal3 s 39200 94120 40000 94240 6 la_data_out[10]
port 460 nsew signal output
rlabel metal3 s 39200 94664 40000 94784 6 la_data_out[11]
port 461 nsew signal output
rlabel metal3 s 39200 95208 40000 95328 6 la_data_out[12]
port 462 nsew signal output
rlabel metal3 s 39200 95752 40000 95872 6 la_data_out[13]
port 463 nsew signal output
rlabel metal3 s 39200 96296 40000 96416 6 la_data_out[14]
port 464 nsew signal output
rlabel metal3 s 39200 96840 40000 96960 6 la_data_out[15]
port 465 nsew signal output
rlabel metal3 s 39200 97384 40000 97504 6 la_data_out[16]
port 466 nsew signal output
rlabel metal3 s 39200 97928 40000 98048 6 la_data_out[17]
port 467 nsew signal output
rlabel metal3 s 39200 98472 40000 98592 6 la_data_out[18]
port 468 nsew signal output
rlabel metal3 s 39200 99016 40000 99136 6 la_data_out[19]
port 469 nsew signal output
rlabel metal3 s 39200 89224 40000 89344 6 la_data_out[1]
port 470 nsew signal output
rlabel metal3 s 39200 99560 40000 99680 6 la_data_out[20]
port 471 nsew signal output
rlabel metal3 s 39200 100104 40000 100224 6 la_data_out[21]
port 472 nsew signal output
rlabel metal3 s 39200 100648 40000 100768 6 la_data_out[22]
port 473 nsew signal output
rlabel metal3 s 39200 101192 40000 101312 6 la_data_out[23]
port 474 nsew signal output
rlabel metal3 s 39200 101736 40000 101856 6 la_data_out[24]
port 475 nsew signal output
rlabel metal3 s 39200 102280 40000 102400 6 la_data_out[25]
port 476 nsew signal output
rlabel metal3 s 39200 102824 40000 102944 6 la_data_out[26]
port 477 nsew signal output
rlabel metal3 s 39200 103368 40000 103488 6 la_data_out[27]
port 478 nsew signal output
rlabel metal3 s 39200 103912 40000 104032 6 la_data_out[28]
port 479 nsew signal output
rlabel metal3 s 39200 104456 40000 104576 6 la_data_out[29]
port 480 nsew signal output
rlabel metal3 s 39200 89768 40000 89888 6 la_data_out[2]
port 481 nsew signal output
rlabel metal3 s 39200 105000 40000 105120 6 la_data_out[30]
port 482 nsew signal output
rlabel metal3 s 39200 105544 40000 105664 6 la_data_out[31]
port 483 nsew signal output
rlabel metal3 s 39200 106088 40000 106208 6 la_data_out[32]
port 484 nsew signal output
rlabel metal3 s 39200 106632 40000 106752 6 la_data_out[33]
port 485 nsew signal output
rlabel metal3 s 39200 107176 40000 107296 6 la_data_out[34]
port 486 nsew signal output
rlabel metal3 s 39200 107720 40000 107840 6 la_data_out[35]
port 487 nsew signal output
rlabel metal3 s 39200 108264 40000 108384 6 la_data_out[36]
port 488 nsew signal output
rlabel metal3 s 39200 108808 40000 108928 6 la_data_out[37]
port 489 nsew signal output
rlabel metal3 s 39200 109352 40000 109472 6 la_data_out[38]
port 490 nsew signal output
rlabel metal3 s 39200 109896 40000 110016 6 la_data_out[39]
port 491 nsew signal output
rlabel metal3 s 39200 90312 40000 90432 6 la_data_out[3]
port 492 nsew signal output
rlabel metal3 s 39200 90856 40000 90976 6 la_data_out[4]
port 493 nsew signal output
rlabel metal3 s 39200 91400 40000 91520 6 la_data_out[5]
port 494 nsew signal output
rlabel metal3 s 39200 91944 40000 92064 6 la_data_out[6]
port 495 nsew signal output
rlabel metal3 s 39200 92488 40000 92608 6 la_data_out[7]
port 496 nsew signal output
rlabel metal3 s 39200 93032 40000 93152 6 la_data_out[8]
port 497 nsew signal output
rlabel metal3 s 39200 93576 40000 93696 6 la_data_out[9]
port 498 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 rst_6502
port 499 nsew signal output
rlabel metal3 s 0 199928 800 200048 6 rst_8x305
port 500 nsew signal output
rlabel metal2 s 37646 219200 37702 220000 6 rst_as1802
port 501 nsew signal output
rlabel metal2 s 36910 219200 36966 220000 6 rst_scrapcpu
port 502 nsew signal output
rlabel metal2 s 9678 219200 9734 220000 6 rst_vliw
port 503 nsew signal output
rlabel metal3 s 39200 130024 40000 130144 6 rst_z80
port 504 nsew signal output
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 505 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 505 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 506 nsew ground bidirectional
rlabel metal3 s 0 50600 800 50720 6 wb_clk_i
port 507 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 wb_rst_i
port 508 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 wbs_ack_o
port 509 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 wbs_adr_i[0]
port 510 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[10]
port 511 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[11]
port 512 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[12]
port 513 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[13]
port 514 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[14]
port 515 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[15]
port 516 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_adr_i[16]
port 517 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[17]
port 518 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[18]
port 519 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[19]
port 520 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[1]
port 521 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[20]
port 522 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[21]
port 523 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[22]
port 524 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[23]
port 525 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[24]
port 526 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[25]
port 527 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[26]
port 528 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[27]
port 529 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_adr_i[28]
port 530 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[29]
port 531 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_adr_i[2]
port 532 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[30]
port 533 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[31]
port 534 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_adr_i[3]
port 535 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[4]
port 536 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[5]
port 537 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[6]
port 538 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[7]
port 539 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[8]
port 540 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_adr_i[9]
port 541 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 wbs_cyc_i
port 542 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 wbs_dat_i[0]
port 543 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 wbs_dat_i[10]
port 544 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 wbs_dat_i[11]
port 545 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 wbs_dat_i[12]
port 546 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 wbs_dat_i[13]
port 547 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wbs_dat_i[14]
port 548 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 wbs_dat_i[15]
port 549 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 wbs_dat_i[16]
port 550 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 wbs_dat_i[17]
port 551 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 wbs_dat_i[18]
port 552 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wbs_dat_i[19]
port 553 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 wbs_dat_i[1]
port 554 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 wbs_dat_i[20]
port 555 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 wbs_dat_i[21]
port 556 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbs_dat_i[22]
port 557 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wbs_dat_i[23]
port 558 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 wbs_dat_i[24]
port 559 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 wbs_dat_i[25]
port 560 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 wbs_dat_i[26]
port 561 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 wbs_dat_i[27]
port 562 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 wbs_dat_i[28]
port 563 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 wbs_dat_i[29]
port 564 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 wbs_dat_i[2]
port 565 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 wbs_dat_i[30]
port 566 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wbs_dat_i[31]
port 567 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 wbs_dat_i[3]
port 568 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 wbs_dat_i[4]
port 569 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 wbs_dat_i[5]
port 570 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 wbs_dat_i[6]
port 571 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 wbs_dat_i[7]
port 572 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 wbs_dat_i[8]
port 573 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 wbs_dat_i[9]
port 574 nsew signal input
rlabel metal3 s 39200 71272 40000 71392 6 wbs_dat_o[0]
port 575 nsew signal output
rlabel metal3 s 39200 76712 40000 76832 6 wbs_dat_o[10]
port 576 nsew signal output
rlabel metal3 s 39200 77256 40000 77376 6 wbs_dat_o[11]
port 577 nsew signal output
rlabel metal3 s 39200 77800 40000 77920 6 wbs_dat_o[12]
port 578 nsew signal output
rlabel metal3 s 39200 78344 40000 78464 6 wbs_dat_o[13]
port 579 nsew signal output
rlabel metal3 s 39200 78888 40000 79008 6 wbs_dat_o[14]
port 580 nsew signal output
rlabel metal3 s 39200 79432 40000 79552 6 wbs_dat_o[15]
port 581 nsew signal output
rlabel metal3 s 39200 79976 40000 80096 6 wbs_dat_o[16]
port 582 nsew signal output
rlabel metal3 s 39200 80520 40000 80640 6 wbs_dat_o[17]
port 583 nsew signal output
rlabel metal3 s 39200 81064 40000 81184 6 wbs_dat_o[18]
port 584 nsew signal output
rlabel metal3 s 39200 81608 40000 81728 6 wbs_dat_o[19]
port 585 nsew signal output
rlabel metal3 s 39200 71816 40000 71936 6 wbs_dat_o[1]
port 586 nsew signal output
rlabel metal3 s 39200 82152 40000 82272 6 wbs_dat_o[20]
port 587 nsew signal output
rlabel metal3 s 39200 82696 40000 82816 6 wbs_dat_o[21]
port 588 nsew signal output
rlabel metal3 s 39200 83240 40000 83360 6 wbs_dat_o[22]
port 589 nsew signal output
rlabel metal3 s 39200 83784 40000 83904 6 wbs_dat_o[23]
port 590 nsew signal output
rlabel metal3 s 39200 84328 40000 84448 6 wbs_dat_o[24]
port 591 nsew signal output
rlabel metal3 s 39200 84872 40000 84992 6 wbs_dat_o[25]
port 592 nsew signal output
rlabel metal3 s 39200 85416 40000 85536 6 wbs_dat_o[26]
port 593 nsew signal output
rlabel metal3 s 39200 85960 40000 86080 6 wbs_dat_o[27]
port 594 nsew signal output
rlabel metal3 s 39200 86504 40000 86624 6 wbs_dat_o[28]
port 595 nsew signal output
rlabel metal3 s 39200 87048 40000 87168 6 wbs_dat_o[29]
port 596 nsew signal output
rlabel metal3 s 39200 72360 40000 72480 6 wbs_dat_o[2]
port 597 nsew signal output
rlabel metal3 s 39200 87592 40000 87712 6 wbs_dat_o[30]
port 598 nsew signal output
rlabel metal3 s 39200 88136 40000 88256 6 wbs_dat_o[31]
port 599 nsew signal output
rlabel metal3 s 39200 72904 40000 73024 6 wbs_dat_o[3]
port 600 nsew signal output
rlabel metal3 s 39200 73448 40000 73568 6 wbs_dat_o[4]
port 601 nsew signal output
rlabel metal3 s 39200 73992 40000 74112 6 wbs_dat_o[5]
port 602 nsew signal output
rlabel metal3 s 39200 74536 40000 74656 6 wbs_dat_o[6]
port 603 nsew signal output
rlabel metal3 s 39200 75080 40000 75200 6 wbs_dat_o[7]
port 604 nsew signal output
rlabel metal3 s 39200 75624 40000 75744 6 wbs_dat_o[8]
port 605 nsew signal output
rlabel metal3 s 39200 76168 40000 76288 6 wbs_dat_o[9]
port 606 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 wbs_stb_i
port 607 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 wbs_we_i
port 608 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 220000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7970844
string GDS_FILE /home/lucah/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/Multiplexer/runs/24_06_04_13_12/results/signoff/multiplexer.magic.gds
string GDS_START 449908
<< end >>

