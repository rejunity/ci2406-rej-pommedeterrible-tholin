* NGSPICE file created from wrapped_8x305.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt wrapped_8x305 custom_settings[0] custom_settings[1] io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27]
+ io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[1]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28]
+ io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst_n vccd1
+ vssd1 wb_clk_i
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3155_ _3842_/Q _3157_/A _3148_/A _3154_/Y vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3086_ _3088_/A _3169_/B _3088_/B vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__or3b_1
X_2106_ _2142_/A _2106_/B vssd1 vssd1 vccd1 vccd1 _2106_/X sky130_fd_sc_hd__or2_1
X_2037_ _2035_/X _2036_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__mux2_1
X_3988_ _4016_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2939_ _2939_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _3201_/B sky130_fd_sc_hd__nor2_1
XANTENNA__2954__A1 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold362 hold743/X vssd1 vssd1 vccd1 vccd1 _1844_/A sky130_fd_sc_hd__buf_1
Xhold351 _3738_/Q vssd1 vssd1 vccd1 vccd1 _2732_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold340 _3865_/Q vssd1 vssd1 vccd1 vccd1 _2407_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _4039_/Q vssd1 vssd1 vccd1 vccd1 _1840_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold395 _3863_/Q vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _3875_/Q vssd1 vssd1 vccd1 vccd1 _3218_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout75_A _1867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output56_A _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3911_ _4101_/CLK _3911_/D vssd1 vssd1 vccd1 vccd1 _3911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3842_ _3846_/CLK _3842_/D vssd1 vssd1 vccd1 vccd1 _3842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3773_ _3794_/CLK _3773_/D vssd1 vssd1 vccd1 vccd1 _3773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2724_ _2720_/A _2723_/X _2735_/S vssd1 vssd1 vccd1 vccd1 _2725_/B sky130_fd_sc_hd__mux2_1
X_2655_ _2345_/X _2573_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2586_ _3720_/Q _2583_/Y _2585_/Y _2579_/Y _2581_/Y vssd1 vssd1 vccd1 vccd1 _2586_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3361__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout105 _2698_/A vssd1 vssd1 vccd1 vccd1 _2805_/A sky130_fd_sc_hd__clkbuf_4
X_3207_ _3693_/Q _3201_/Y _3206_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__o211a_1
X_3138_ _3138_/A _3138_/B vssd1 vssd1 vccd1 vccd1 _3138_/Y sky130_fd_sc_hd__nor2_1
X_3069_ _3832_/Q _2923_/B _2922_/Y _2935_/B vssd1 vssd1 vccd1 vccd1 _3069_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold170 _3390_/X vssd1 vssd1 vccd1 vccd1 _3954_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _3402_/X vssd1 vssd1 vccd1 vccd1 _3964_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _3702_/Q vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2538__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1969__A2 _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2091__B2 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2034__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _3970_/Q _4067_/Q _4059_/Q _4051_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2441_/B sky130_fd_sc_hd__mux4_1
XANTENNA__3343__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2371_ _2376_/A _2376_/C vssd1 vssd1 vccd1 vccd1 _2484_/B sky130_fd_sc_hd__nand2_1
X_4110_ _4113_/CLK _4110_/D vssd1 vssd1 vccd1 vccd1 _4110_/Q sky130_fd_sc_hd__dfxtp_1
X_4041_ _4092_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _4041_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2082__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3825_ _3846_/CLK _3825_/D vssd1 vssd1 vccd1 vccd1 _3825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3756_ _3803_/CLK _3756_/D vssd1 vssd1 vccd1 vccd1 _3756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2707_ _2678_/X _2690_/Y _2706_/X vssd1 vssd1 vccd1 vccd1 _3728_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3687_ hold609/X _2681_/Y _2688_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3687_/X sky130_fd_sc_hd__o211a_1
X_2638_ _2637_/B _2637_/C hold1/X vssd1 vssd1 vccd1 vccd1 _2638_/Y sky130_fd_sc_hd__a21oi_1
X_2569_ hold520/X _2556_/Y _2568_/X _2555_/X _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3694_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2119__S _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3325__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1940_ _2616_/A _2616_/B _2616_/C vssd1 vssd1 vccd1 vccd1 _1942_/B sky130_fd_sc_hd__and3_2
XANTENNA__2064__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1871_ _2923_/B vssd1 vssd1 vccd1 vccd1 _3123_/B sky130_fd_sc_hd__inv_2
X_3610_ _3637_/A0 hold23/X _3612_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3541_ _3529_/A _3525_/B _3528_/B vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3472_ _3472_/A _3496_/S vssd1 vssd1 vccd1 vccd1 _3472_/Y sky130_fd_sc_hd__nand2_1
X_2423_ _2422_/X _2420_/Y _2484_/A vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__mux2_1
X_2354_ _2737_/C _2351_/X _2352_/X _2353_/Y vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__o22a_1
X_2285_ _2285_/A _2285_/B _2284_/X vssd1 vssd1 vccd1 vccd1 _2285_/X sky130_fd_sc_hd__or3b_1
X_4024_ _4031_/CLK _4024_/D vssd1 vssd1 vccd1 vccd1 _4024_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3252__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _4092_/CLK _3808_/D vssd1 vssd1 vccd1 vccd1 _3808_/Q sky130_fd_sc_hd__dfxtp_2
X_3739_ _3803_/CLK _3739_/D vssd1 vssd1 vccd1 vccd1 _3739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2046__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2506__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _2068_/X _2069_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2972_ _3199_/A _3817_/Q vssd1 vssd1 vccd1 vccd1 _2972_/Y sky130_fd_sc_hd__nand2_1
X_1923_ _2230_/A _3507_/A _2376_/A _2369_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _3322_/A
+ sky130_fd_sc_hd__o2111a_4
XFILLER_0_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1854_ _1854_/A vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3537__A1 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold703 _3070_/Y vssd1 vssd1 vccd1 vccd1 _3071_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3524_ _1846_/A _3564_/B _3522_/Y _3523_/X _3587_/A vssd1 vssd1 vccd1 vccd1 _4032_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold725 _3836_/Q vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _3829_/Q vssd1 vssd1 vccd1 vccd1 _3060_/B sky130_fd_sc_hd__clkbuf_2
Xhold736 _4097_/Q vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
X_3455_ _3455_/A _3675_/B vssd1 vssd1 vccd1 vccd1 _3470_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold747 _3707_/Q vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
X_2406_ _1887_/Y _2405_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2406_/X sky130_fd_sc_hd__mux2_1
X_3386_ _3454_/A _3631_/B vssd1 vssd1 vccd1 vccd1 _3604_/C sky130_fd_sc_hd__or2_1
X_2337_ _2508_/A _2337_/B vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2268_ _2268_/A _2315_/B _2327_/B vssd1 vssd1 vccd1 vccd1 _2376_/B sky130_fd_sc_hd__and3_1
X_4007_ _4011_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
X_2199_ _2378_/A _2378_/B vssd1 vssd1 vccd1 vccd1 _2424_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4088_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3519__A1 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3519__B2 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2042__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _2531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _1840_/Y _1855_/Y _3496_/S vssd1 vssd1 vccd1 vccd1 _3240_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3812__D _3812_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3171_ _3171_/A _3294_/B vssd1 vssd1 vccd1 vccd1 _3189_/S sky130_fd_sc_hd__nand2_8
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2120_/X _2121_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2122_/X sky130_fd_sc_hd__mux2_1
X_2053_ _3767_/Q _3751_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2053_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2955_ hold643/X _2940_/X _3114_/A vssd1 vssd1 vccd1 vccd1 _2955_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2886_ _2674_/X _2871_/X _2885_/X vssd1 vssd1 vccd1 vccd1 _3802_/D sky130_fd_sc_hd__a21o_1
X_1906_ _1906_/A _2180_/B vssd1 vssd1 vccd1 vccd1 _2646_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold500 _2944_/Y vssd1 vssd1 vccd1 vccd1 _3810_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _3923_/Q vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _3814_/Q vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _3921_/Q vssd1 vssd1 vccd1 vccd1 _3324_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold533 _2800_/X vssd1 vssd1 vccd1 vccd1 _3764_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3507_/A _3507_/B vssd1 vssd1 vccd1 vccd1 _3507_/X sky130_fd_sc_hd__and2_1
Xhold588 _3246_/X vssd1 vssd1 vccd1 vccd1 _3247_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold577 _3826_/Q vssd1 vssd1 vccd1 vccd1 _3120_/A sky130_fd_sc_hd__buf_2
Xhold566 _3668_/X vssd1 vssd1 vccd1 vccd1 _4099_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _3912_/Q vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3438_ _3633_/A0 hold121/X _3444_/S vssd1 vssd1 vccd1 vccd1 _3438_/X sky130_fd_sc_hd__mux2_1
Xhold599 _3828_/Q vssd1 vssd1 vccd1 vccd1 _2990_/D sky130_fd_sc_hd__clkbuf_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _2667_/X _3358_/X _3368_/X vssd1 vssd1 vccd1 vccd1 _3941_/D sky130_fd_sc_hd__a21o_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput31 _2592_/C vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
Xoutput42 _3836_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
Xoutput53 _3635_/A0 vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__2037__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2740_ _2738_/X _2739_/X _2740_/S vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2671_ _2462_/X _2677_/B _2670_/Y vssd1 vssd1 vccd1 vccd1 _2671_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_78_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2479__A1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3676__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3223_ _3458_/A _2681_/Y _3222_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3223_/X sky130_fd_sc_hd__o211a_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _3157_/A _3154_/B vssd1 vssd1 vccd1 vccd1 _3154_/Y sky130_fd_sc_hd__nor2_1
X_3085_ _3099_/C _3125_/A vssd1 vssd1 vccd1 vccd1 _3088_/B sky130_fd_sc_hd__or2_1
XANTENNA__2736__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2105_ _3716_/Q _3728_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2106_/B sky130_fd_sc_hd__mux2_1
X_2036_ _3772_/Q _3788_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2036_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _4011_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2938_ _3658_/A _2936_/X _3494_/S _3601_/A vssd1 vssd1 vccd1 vccd1 _3808_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2954__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2869_ _2869_/A _2869_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__and3_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold352 _2625_/Y vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _4096_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _3207_/X vssd1 vssd1 vccd1 vccd1 _3865_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold363 _3232_/X vssd1 vssd1 vccd1 vccd1 _3233_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _3240_/X vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _3203_/X vssd1 vssd1 vccd1 vccd1 _3863_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _3219_/X vssd1 vssd1 vccd1 vccd1 _3875_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3667__A0 _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout68_A _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3419__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A _3467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2945__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3910_ _4105_/CLK _3910_/D vssd1 vssd1 vccd1 vccd1 _3910_/Q sky130_fd_sc_hd__dfxtp_1
X_3841_ _3846_/CLK _3841_/D vssd1 vssd1 vccd1 vccd1 _3841_/Q sky130_fd_sc_hd__dfxtp_1
X_3772_ _3795_/CLK _3772_/D vssd1 vssd1 vccd1 vccd1 _3772_/Q sky130_fd_sc_hd__dfxtp_1
X_2723_ _2327_/B _2721_/X _2734_/S vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__mux2_1
X_2654_ _2869_/A _2654_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__and3_1
X_2585_ _2585_/A _2585_/B vssd1 vssd1 vccd1 vccd1 _2585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout106 _2698_/A vssd1 vssd1 vccd1 vccd1 _2863_/A sky130_fd_sc_hd__clkbuf_2
X_3206_ _1889_/Y _3201_/A _2410_/B _2407_/B vssd1 vssd1 vccd1 vccd1 _3206_/X sky130_fd_sc_hd__a31o_1
X_3137_ _2988_/B _3133_/B _3134_/Y _3120_/D vssd1 vssd1 vccd1 vccd1 _3138_/B sky130_fd_sc_hd__o2bb2a_1
X_3068_ _3065_/B _3057_/X _3067_/X hold710/X _3497_/A vssd1 vssd1 vccd1 vccd1 _3068_/X
+ sky130_fd_sc_hd__o311a_1
X_2019_ _2015_/X _2018_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold160 _3419_/X vssd1 vssd1 vccd1 vccd1 _3978_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2140__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 _4111_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold193 _4057_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _2602_/X vssd1 vssd1 vccd1 vccd1 _3702_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1969__A3 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ _2376_/A _2376_/C vssd1 vssd1 vccd1 vccd1 _2373_/B sky130_fd_sc_hd__and2_1
X_4040_ _4045_/CLK _4040_/D vssd1 vssd1 vccd1 vccd1 _4040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3824_ _3862_/CLK _3824_/D vssd1 vssd1 vccd1 vccd1 _3824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_46_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3755_ _3795_/CLK _3755_/D vssd1 vssd1 vccd1 vccd1 _3755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2706_ _2813_/A _2706_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2706_/X sky130_fd_sc_hd__and3_1
X_3686_ hold688/X _2681_/Y _2686_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3686_/X sky130_fd_sc_hd__o211a_1
X_2637_ hold1/X _2637_/B _2637_/C vssd1 vssd1 vccd1 vccd1 _2642_/B sky130_fd_sc_hd__and3_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2568_ _2393_/B _2567_/X _2556_/Y vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__a21bo_1
X_2499_ _2564_/A _2499_/B vssd1 vssd1 vccd1 vccd1 _2499_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3270__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1870_ _2935_/B vssd1 vssd1 vccd1 vccd1 _3275_/B sky130_fd_sc_hd__inv_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3540_ _3540_/A _3540_/B vssd1 vssd1 vccd1 vccd1 _3543_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3471_ hold282/X _3470_/B _3470_/Y _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3471_/X sky130_fd_sc_hd__o211a_1
X_2422_ _2378_/A _2424_/A _2424_/C _2424_/B vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__a31o_1
X_2353_ _2352_/A _2352_/B _2737_/C vssd1 vssd1 vccd1 vccd1 _2353_/Y sky130_fd_sc_hd__o21ai_1
X_2284_ _2260_/X _2283_/X _2247_/X vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__a21o_1
X_4023_ _4092_/CLK _4023_/D vssd1 vssd1 vccd1 vccd1 _4023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2744__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3807_ _4095_/CLK _3807_/D vssd1 vssd1 vccd1 vccd1 _3807_/Q sky130_fd_sc_hd__dfxtp_1
X_1999_ _1987_/A _1998_/X _3554_/B _1918_/X vssd1 vssd1 vccd1 vccd1 _2192_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3738_ _3803_/CLK _3738_/D vssd1 vssd1 vccd1 vccd1 _3738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3669_ _2119_/S hold592/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2818__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output31_A _2592_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ _3157_/A _3081_/A _2957_/Y vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ _2230_/A _3507_/A _2376_/A vssd1 vssd1 vccd1 vccd1 _2834_/B sky130_fd_sc_hd__o21ai_2
X_1853_ _1853_/A vssd1 vssd1 vccd1 vccd1 _1853_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 _4037_/Q vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 _3887_/Q vssd1 vssd1 vccd1 vccd1 _1854_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ _2619_/A _3554_/B hold368/X vssd1 vssd1 vccd1 vccd1 _3523_/X sky130_fd_sc_hd__a21o_1
Xhold726 _3113_/X vssd1 vssd1 vccd1 vccd1 _3114_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 _3739_/Q vssd1 vssd1 vccd1 vccd1 _2738_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3454_ _3454_/A _3872_/Q _3871_/Q vssd1 vssd1 vccd1 vccd1 _3675_/B sky130_fd_sc_hd__or3b_4
X_2405_ _3720_/Q _2402_/Y _2404_/Y _2398_/Y _2400_/Y vssd1 vssd1 vccd1 vccd1 _2405_/X
+ sky130_fd_sc_hd__a32o_1
X_3385_ _3872_/Q _3871_/Q vssd1 vssd1 vccd1 vccd1 _3631_/B sky130_fd_sc_hd__nand2_1
X_2336_ _2334_/Y _2335_/X _2571_/B vssd1 vssd1 vccd1 vccd1 _2337_/B sky130_fd_sc_hd__a21oi_1
X_2267_ _2227_/S _3502_/B _3554_/A vssd1 vssd1 vccd1 vccd1 _2267_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4006_ _4014_/CLK _4006_/D vssd1 vssd1 vccd1 vccd1 _4006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2198_ _2421_/A _2327_/B vssd1 vssd1 vccd1 vccd1 _2424_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_A input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3216__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_6 _1862_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3171_/A _3294_/B vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__and2_1
X_2121_ _3934_/Q _3926_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2121_/X sky130_fd_sc_hd__mux2_1
X_2052_ _2050_/X _2051_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3207__A1 _3693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2954_ _3633_/A0 _2940_/X _2953_/Y vssd1 vssd1 vccd1 vccd1 _3815_/D sky130_fd_sc_hd__a21oi_1
X_2885_ _2887_/A _2885_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__and3_1
X_1905_ _1987_/A _2616_/C vssd1 vssd1 vccd1 vccd1 _2269_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold501 _3709_/Q vssd1 vssd1 vccd1 vccd1 _2654_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _3809_/Q vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3391__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 _3325_/X vssd1 vssd1 vccd1 vccd1 _3921_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold534 _3788_/Q vssd1 vssd1 vccd1 vccd1 _2855_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3506_/A _3506_/B vssd1 vssd1 vccd1 vccd1 _3506_/X sky130_fd_sc_hd__xor2_2
Xhold545 _3872_/Q vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout100_A _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 _3821_/Q vssd1 vssd1 vccd1 vccd1 _2891_/A sky130_fd_sc_hd__buf_1
Xhold578 _3000_/Y vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _3290_/X vssd1 vssd1 vccd1 vccd1 _3291_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ _1861_/Y hold231/X _3444_/S vssd1 vssd1 vccd1 vccd1 _3437_/X sky130_fd_sc_hd__mux2_1
Xhold589 hold736/X vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3654_/A _3368_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3368_/X sky130_fd_sc_hd__and3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _3321_/A _2296_/X _2297_/X _2093_/B vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__o22a_1
X_3299_ input6/X hold611/X _3301_/S vssd1 vssd1 vccd1 vccd1 _3299_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2932__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2143__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3382__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput43 _3809_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_12
Xoutput32 _2939_/B vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
Xoutput54 _3636_/A0 vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ _2670_/A _2677_/B vssd1 vssd1 vccd1 vccd1 _2670_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2053__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3222_ _3222_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _3222_/X sky130_fd_sc_hd__or2_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _3163_/A _2961_/X _3157_/B vssd1 vssd1 vccd1 vccd1 _3154_/B sky130_fd_sc_hd__a21oi_1
X_2104_ _2102_/X _2103_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2104_/X sky130_fd_sc_hd__mux2_1
X_3084_ _3125_/A vssd1 vssd1 vccd1 vccd1 _3084_/Y sky130_fd_sc_hd__inv_2
X_2035_ _3764_/Q _3748_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3986_ _4016_/CLK _3986_/D vssd1 vssd1 vccd1 vccd1 _3986_/Q sky130_fd_sc_hd__dfxtp_1
X_2937_ _2937_/A _3065_/B vssd1 vssd1 vccd1 vccd1 _2937_/X sky130_fd_sc_hd__or2_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2868_ _2674_/X _2853_/X _2867_/X vssd1 vssd1 vccd1 vccd1 _3794_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold320 hold733/X vssd1 vssd1 vccd1 vccd1 _2630_/A sky130_fd_sc_hd__buf_1
X_2799_ _2813_/A _2799_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2799_/X sky130_fd_sc_hd__and3_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 hold734/X vssd1 vssd1 vccd1 vccd1 _2624_/A sky130_fd_sc_hd__buf_1
Xhold353 _2626_/X vssd1 vssd1 vccd1 vccd1 _2627_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _3665_/X vssd1 vssd1 vccd1 vccd1 _4096_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _3932_/Q vssd1 vssd1 vccd1 vccd1 _3348_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _3747_/Q vssd1 vssd1 vccd1 vccd1 _2758_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _3866_/Q vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 _3790_/Q vssd1 vssd1 vccd1 vccd1 _2859_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2330__A1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2330__B2 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _3846_/CLK _3840_/D vssd1 vssd1 vccd1 vccd1 _3840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3771_ _3795_/CLK _3771_/D vssd1 vssd1 vccd1 vccd1 _3771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2722_ _3554_/A _2733_/S _2615_/B vssd1 vssd1 vccd1 vccd1 _2735_/S sky130_fd_sc_hd__a21oi_2
X_2653_ _3341_/A _3258_/A vssd1 vssd1 vccd1 vccd1 _2676_/C sky130_fd_sc_hd__or2_2
X_2584_ hold99/A _3897_/Q _3703_/Q hold39/A _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2585_/B sky130_fd_sc_hd__mux4_2
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout107 _2813_/A vssd1 vssd1 vccd1 vccd1 _2869_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3649__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3205_ hold730/X _3201_/Y _3204_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__o211a_1
X_3136_ _3136_/A _3136_/B _3136_/C vssd1 vssd1 vccd1 vccd1 _3138_/A sky130_fd_sc_hd__or3_1
X_3067_ _3123_/A _3067_/B vssd1 vssd1 vccd1 vccd1 _3067_/X sky130_fd_sc_hd__xor2_1
X_2018_ _2016_/X _2017_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2018_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ _4073_/CLK _3969_/D vssd1 vssd1 vccd1 vccd1 _3969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold161 _4052_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold150 _3619_/X vssd1 vssd1 vccd1 vccd1 _4063_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _3612_/X vssd1 vssd1 vccd1 vccd1 _4057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _3681_/X vssd1 vssd1 vccd1 vccd1 _4111_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _4061_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout80_A _1862_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3823_ _4077_/CLK _3823_/D vssd1 vssd1 vccd1 vccd1 _3823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4016_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _3794_/CLK _3754_/D vssd1 vssd1 vccd1 vccd1 _3754_/Q sky130_fd_sc_hd__dfxtp_1
X_2705_ _2674_/X _2690_/Y _2704_/X vssd1 vssd1 vccd1 vccd1 _3727_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3685_ hold520/X _2681_/Y _2684_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3685_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2790__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2636_ _2637_/B _2640_/B _2635_/Y _3227_/A vssd1 vssd1 vccd1 vccd1 _3706_/D sky130_fd_sc_hd__o211a_1
X_2567_ _2566_/X input9/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2498_ hold41/A _4109_/Q _3964_/Q hold97/A _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2499_/B sky130_fd_sc_hd__mux4_1
X_3119_ _3120_/A _3119_/B _3120_/D vssd1 vssd1 vccd1 vccd1 _3308_/A sky130_fd_sc_hd__or3_1
X_4099_ _4101_/CLK _4099_/D vssd1 vssd1 vccd1 vccd1 _4099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3007__C1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2151__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2297__B1 _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2772__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3470_ _3695_/Q _3470_/B vssd1 vssd1 vccd1 vccd1 _3470_/Y sky130_fd_sc_hd__nand2_1
X_2421_ _2421_/A _2484_/B vssd1 vssd1 vccd1 vccd1 _2424_/C sky130_fd_sc_hd__nand2_1
X_2352_ _2352_/A _2352_/B vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__and2_1
XFILLER_0_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2283_ _2345_/S _2338_/B _2350_/B _2272_/Y vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__a211o_1
X_4022_ _4031_/CLK _4022_/D vssd1 vssd1 vccd1 vccd1 _4022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3806_ _4105_/CLK _3806_/D vssd1 vssd1 vccd1 vccd1 _3806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3575__B _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3737_ _4101_/CLK _3737_/D vssd1 vssd1 vccd1 vccd1 _3737_/Q sky130_fd_sc_hd__dfxtp_1
X_1998_ _1918_/X _1997_/X _3544_/S vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3668_ _2151_/S hold565/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__mux2_1
X_2619_ _2619_/A _2619_/B _3584_/A vssd1 vssd1 vccd1 vccd1 _3592_/B sky130_fd_sc_hd__and3_2
X_3599_ _2621_/A _2613_/Y _3596_/Y _3598_/X _2887_/A vssd1 vssd1 vccd1 vccd1 _3599_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2056__S _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output24_A _1976_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2970_ _3163_/A _3134_/C _3075_/B _2968_/B _3150_/B vssd1 vssd1 vccd1 vccd1 _3081_/A
+ sky130_fd_sc_hd__a311o_1
X_1921_ _2230_/A _3507_/A _2376_/A vssd1 vssd1 vccd1 vccd1 _2710_/B sky130_fd_sc_hd__o21a_2
X_1852_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2745__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3522_ _3554_/B _3522_/B vssd1 vssd1 vccd1 vccd1 _3522_/Y sky130_fd_sc_hd__nor2_1
Xhold716 _2912_/X vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold705 _3834_/Q vssd1 vssd1 vccd1 vccd1 _3275_/A sky130_fd_sc_hd__clkbuf_2
Xhold727 _3830_/Q vssd1 vssd1 vccd1 vccd1 _3036_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3453_ _3639_/A0 hold69/X _3453_/S vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__mux2_1
Xhold738 _4040_/Q vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
X_2404_ _2564_/A _2404_/B vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__nand2_1
X_3384_ _3639_/A0 hold99/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__mux2_1
X_2335_ _2362_/S _2670_/A _2328_/Y _2347_/S vssd1 vssd1 vccd1 vccd1 _2335_/X sky130_fd_sc_hd__a211o_1
X_2266_ _2279_/S _2266_/B _2266_/C vssd1 vssd1 vccd1 vccd1 _2266_/X sky130_fd_sc_hd__or3_1
X_4005_ _4016_/CLK _4005_/D vssd1 vssd1 vccd1 vccd1 _4005_/Q sky130_fd_sc_hd__dfxtp_1
X_2197_ _2197_/A _2197_/B vssd1 vssd1 vccd1 vccd1 _2197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _3965_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _4087_/Q _3942_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2120_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3794_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2051_ _3743_/Q _3759_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2051_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1910__C _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2953_ hold598/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2953_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1904_ _4104_/Q _1890_/Y _1902_/X vssd1 vssd1 vccd1 vccd1 _2616_/C sky130_fd_sc_hd__o21ai_4
X_2884_ _2671_/X _2871_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _3801_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2718__B2 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 _2656_/X vssd1 vssd1 vccd1 vccd1 _3709_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _2942_/Y vssd1 vssd1 vccd1 vccd1 _3809_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold535 _2856_/X vssd1 vssd1 vccd1 vccd1 _3788_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3505_/A _3505_/B vssd1 vssd1 vccd1 vccd1 _3505_/X sky130_fd_sc_hd__or2_1
Xhold524 _3900_/Q vssd1 vssd1 vccd1 vccd1 _3263_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _2987_/X vssd1 vssd1 vccd1 vccd1 _3821_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _3002_/Y vssd1 vssd1 vccd1 vccd1 _3826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _3910_/Q vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _2685_/X vssd1 vssd1 vccd1 vccd1 _3718_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3436_ _3613_/C _3455_/A vssd1 vssd1 vccd1 vccd1 _3444_/S sky130_fd_sc_hd__or2_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _2664_/X _3358_/X _3366_/X vssd1 vssd1 vccd1 vccd1 _3940_/D sky130_fd_sc_hd__a21o_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2295_/X _2571_/A _2301_/Y _2304_/Y _2317_/Y vssd1 vssd1 vccd1 vccd1 _2318_/X
+ sky130_fd_sc_hd__a311o_1
X_3298_ _3601_/A _3298_/B vssd1 vssd1 vccd1 vccd1 _3915_/D sky130_fd_sc_hd__and2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2249_ _2222_/B _2187_/X _2194_/A vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2590__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput33 _1944_/X vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
XANTENNA__1932__A2 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput44 _3810_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput55 _3637_/A0 vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2948__A1 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3373__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1923__A2 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2559__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3221_ _3460_/A _2681_/Y _3220_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__o211a_1
X_3152_ hold296/X _3165_/B _3151_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__o211a_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _3936_/Q _3928_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2103_/X sky130_fd_sc_hd__mux2_1
X_3083_ _3834_/Q _3833_/Q _3829_/Q _3830_/Q vssd1 vssd1 vccd1 vccd1 _3125_/A sky130_fd_sc_hd__or4b_2
X_2034_ _2032_/X _2033_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2034_/X sky130_fd_sc_hd__mux2_1
X_3985_ _4016_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2936_ _3065_/B _3073_/A vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__and2b_1
X_2867_ _2869_/A _2867_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__and3_1
XFILLER_0_60_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold310 _3819_/Q vssd1 vssd1 vccd1 vccd1 _2984_/B sky130_fd_sc_hd__clkdlybuf4s25_1
X_2798_ _3340_/A _2854_/A vssd1 vssd1 vccd1 vccd1 _2813_/C sky130_fd_sc_hd__nand2_2
Xhold321 _3574_/X vssd1 vssd1 vccd1 vccd1 _4039_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold738/X vssd1 vssd1 vccd1 vccd1 _3575_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold343 _2629_/B vssd1 vssd1 vccd1 vccd1 _2630_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold387 _2759_/X vssd1 vssd1 vccd1 vccd1 _3747_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _3209_/X vssd1 vssd1 vccd1 vccd1 _3866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _3864_/Q vssd1 vssd1 vccd1 vccd1 _2407_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _3878_/Q vssd1 vssd1 vccd1 vccd1 _3224_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ _3633_/A0 hold159/X _3425_/S vssd1 vssd1 vccd1 vccd1 _3419_/X sky130_fd_sc_hd__mux2_1
Xhold398 _3929_/Q vssd1 vssd1 vccd1 vccd1 _3342_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2646__C _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2154__S _2160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1993__S _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3355__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3770_ _3794_/CLK _3770_/D vssd1 vssd1 vccd1 vccd1 _3770_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3594__A1 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2721_ _2720_/Y _3551_/B _2733_/S vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2652_ _3341_/A _3258_/A vssd1 vssd1 vccd1 vccd1 _2652_/Y sky130_fd_sc_hd__nor2_2
X_2583_ _2585_/A _2583_/B vssd1 vssd1 vccd1 vccd1 _2583_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout108 _2698_/A vssd1 vssd1 vccd1 vccd1 _2813_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3204_ _1889_/Y _3201_/A _2410_/B _2407_/C vssd1 vssd1 vccd1 vccd1 _3204_/X sky130_fd_sc_hd__a31o_1
X_3135_ _3120_/D _3134_/Y _3121_/B vssd1 vssd1 vccd1 vccd1 _3136_/C sky130_fd_sc_hd__o21a_1
X_3066_ _3123_/B _3276_/A vssd1 vssd1 vccd1 vccd1 _3067_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2017_ _3773_/Q _3789_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2763__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2085__A1 _3693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3968_ _4113_/CLK _3968_/D vssd1 vssd1 vccd1 vccd1 _3968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2919_ _2919_/A _2919_/B vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3585__B2 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3899_ _3902_/CLK _3899_/D vssd1 vssd1 vccd1 vccd1 _3899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3337__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold162 _3607_/X vssd1 vssd1 vccd1 vccd1 _4052_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 _3634_/X vssd1 vssd1 vccd1 vccd1 _4076_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _4051_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _3968_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _3617_/X vssd1 vssd1 vccd1 vccd1 _4061_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _4001_/Q vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2673__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2392__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2000__A1 _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2059__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2067__A1 _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3822_ _4077_/CLK _3822_/D vssd1 vssd1 vccd1 vccd1 _3822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3753_ _3794_/CLK _3753_/D vssd1 vssd1 vccd1 vccd1 _3753_/Q sky130_fd_sc_hd__dfxtp_1
X_2704_ _2813_/A _2704_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2704_/X sky130_fd_sc_hd__and3_1
X_3684_ hold559/X _2681_/Y _2682_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3684_/X sky130_fd_sc_hd__o211a_1
X_2635_ _1959_/C _2734_/S _3589_/A _2634_/Y _2640_/B vssd1 vssd1 vccd1 vccd1 _2635_/Y
+ sky130_fd_sc_hd__o221ai_1
XANTENNA__2527__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2566_ _1881_/Y _2565_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2758__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2497_ _2564_/A _2496_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2497_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3118_ _3828_/Q _3118_/B _3140_/B _3140_/C vssd1 vssd1 vccd1 vccd1 _3121_/B sky130_fd_sc_hd__or4_1
X_4098_ _4105_/CLK _4098_/D vssd1 vssd1 vccd1 vccd1 _4098_/Q sky130_fd_sc_hd__dfxtp_1
X_3049_ _3861_/Q _3050_/C _3050_/A vssd1 vssd1 vccd1 vccd1 _3049_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3255__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2297__A1 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3549__A1 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout90 _3717_/Q vssd1 vssd1 vccd1 vccd1 _2584_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2420_ _2420_/A vssd1 vssd1 vccd1 vccd1 _2420_/Y sky130_fd_sc_hd__inv_2
X_2351_ _1945_/Y _2350_/B _2352_/B _2181_/A vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__a2bb2o_1
X_2282_ _2345_/S _2338_/B _2272_/Y vssd1 vssd1 vccd1 vccd1 _2352_/A sky130_fd_sc_hd__a21oi_1
X_4021_ _4029_/CLK _4021_/D vssd1 vssd1 vccd1 vccd1 _4021_/Q sky130_fd_sc_hd__dfxtp_1
X_3805_ _4095_/CLK _3805_/D vssd1 vssd1 vccd1 vccd1 _3805_/Q sky130_fd_sc_hd__dfxtp_1
X_1997_ _2327_/B _3581_/A _2227_/S vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3736_ _4101_/CLK _3736_/D vssd1 vssd1 vccd1 vccd1 _3736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3667_ _2153_/S hold286/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__mux2_1
X_2618_ _3589_/A vssd1 vssd1 vccd1 vccd1 _3596_/B sky130_fd_sc_hd__inv_2
X_3598_ _3596_/B _2720_/B _3597_/X _2615_/B vssd1 vssd1 vccd1 vccd1 _3598_/X sky130_fd_sc_hd__a31o_1
X_2549_ _2570_/A _2549_/B vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2670__B _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3400__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1920_ _1987_/A _2616_/C _2153_/S vssd1 vssd1 vccd1 vccd1 _2376_/A sky130_fd_sc_hd__or3_2
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1851_ _3906_/Q vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__inv_2
X_3521_ _3517_/Y _3520_/Y _3544_/S vssd1 vssd1 vccd1 vccd1 _3522_/B sky130_fd_sc_hd__mux2_1
Xhold728 _4010_/Q vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 _3008_/B vssd1 vssd1 vccd1 vccd1 _3073_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _3065_/B vssd1 vssd1 vccd1 vccd1 _3009_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _1867_/Y hold5/X _3453_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
Xhold739 _3862_/Q vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
X_2403_ _3945_/Q hold73/A _3696_/Q _4074_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2404_/B sky130_fd_sc_hd__mux4_1
X_3383_ _3682_/A0 hold83/X _3384_/S vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
X_2334_ _2349_/B _2332_/X _2347_/S _3540_/A vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__o211ai_1
X_2265_ _2263_/X _2264_/X _2238_/B vssd1 vssd1 vccd1 vccd1 _2266_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__1940__A _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _4016_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
X_2196_ _2093_/B _2191_/X _2195_/X _2094_/Y vssd1 vssd1 vccd1 vccd1 _2197_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2433__A1 _3458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3630__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _4014_/CLK _3719_/D vssd1 vssd1 vccd1 vccd1 _3719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3621__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 _3809_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ hold31/A _3799_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2952_ _3634_/A0 _2940_/X _2951_/Y vssd1 vssd1 vccd1 vccd1 _3814_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__3612__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1903_ hold639/X _1890_/Y _1902_/X vssd1 vssd1 vccd1 vccd1 _2180_/B sky130_fd_sc_hd__o21a_4
X_2883_ _2887_/A _2883_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold536 _3812_/Q vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold514 _3753_/Q vssd1 vssd1 vccd1 vccd1 _2773_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _3748_/Q vssd1 vssd1 vccd1 vccd1 _2763_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3504_ _3507_/A _2277_/B _3502_/X _3554_/A vssd1 vssd1 vccd1 vccd1 _3505_/B sky130_fd_sc_hd__a31o_1
Xhold503 _3785_/Q vssd1 vssd1 vccd1 vccd1 _2847_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _3639_/A0 hold81/X _3435_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
Xhold547 _3813_/Q vssd1 vssd1 vccd1 vccd1 hold547/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold558 _3286_/X vssd1 vssd1 vccd1 vccd1 _3287_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _3871_/Q vssd1 vssd1 vccd1 vccd1 _2682_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _3654_/A _3366_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3366_/X sky130_fd_sc_hd__and3_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2314_/X _2316_/X _2571_/A vssd1 vssd1 vccd1 vccd1 _2317_/Y sky130_fd_sc_hd__a21oi_1
X_3297_ input5/X hold625/X _3301_/S vssd1 vssd1 vccd1 vccd1 _3297_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2248_ _2222_/C _2221_/C _1995_/Y vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2179_ _2177_/Y _2179_/B vssd1 vssd1 vccd1 vccd1 _2291_/A sky130_fd_sc_hd__and2b_1
XANTENNA__3603__B1 _3467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput34 _2940_/A vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
Xoutput45 _3811_/Q vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_12
Xoutput56 _3682_/A0 vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XANTENNA__2676__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2948__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2559__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ _3876_/Q _3224_/B vssd1 vssd1 vccd1 vccd1 _3220_/X sky130_fd_sc_hd__or2_1
XANTENNA__2333__B1 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3151_ hold288/X _3157_/A _3148_/A _3150_/Y vssd1 vssd1 vccd1 vccd1 _3151_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2884__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2102_ _4089_/Q _3944_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__mux2_1
X_3082_ _2988_/B _3169_/B _3157_/A vssd1 vssd1 vccd1 vccd1 _3136_/A sky130_fd_sc_hd__a21o_1
X_2033_ _3740_/Q _3756_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2033_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2525__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3984_ _4113_/CLK hold96/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2935_ _3099_/A _2935_/B _3132_/A vssd1 vssd1 vccd1 vccd1 _3008_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2866_ _2671_/X _2853_/X _2865_/X vssd1 vssd1 vccd1 vccd1 _3793_/D sky130_fd_sc_hd__a21o_1
Xhold311 _2980_/X vssd1 vssd1 vccd1 vccd1 _3819_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold300 _3805_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
X_2797_ _3340_/A _2854_/A vssd1 vssd1 vccd1 vccd1 _2797_/X sky130_fd_sc_hd__and2_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold333 _3242_/X vssd1 vssd1 vccd1 vccd1 _3243_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _2631_/X vssd1 vssd1 vccd1 vccd1 _2632_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 _3831_/Q vssd1 vssd1 vccd1 vccd1 _2923_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2572__A0 hold559/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 _3716_/Q vssd1 vssd1 vccd1 vccd1 _2676_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _3205_/X vssd1 vssd1 vccd1 vccd1 _3864_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _3225_/X vssd1 vssd1 vccd1 vccd1 _3878_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 _3343_/X vssd1 vssd1 vccd1 vccd1 _3929_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ _3676_/A0 hold105/X _3425_/S vssd1 vssd1 vccd1 vccd1 _3418_/X sky130_fd_sc_hd__mux2_1
Xhold388 _3802_/Q vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3349_ _2664_/X _3340_/X _3348_/X vssd1 vssd1 vccd1 vccd1 _3932_/D sky130_fd_sc_hd__a21o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2646__D _2646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2866__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2720_ _2720_/A _2720_/B vssd1 vssd1 vccd1 vccd1 _2720_/Y sky130_fd_sc_hd__xnor2_1
X_2651_ _3321_/B _3641_/A _3321_/A vssd1 vssd1 vccd1 vccd1 _3258_/A sky130_fd_sc_hd__or3b_4
XANTENNA__2080__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2582_ hold95/A _4113_/Q _3968_/Q _3960_/Q _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2583_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout109 _3656_/A vssd1 vssd1 vccd1 vccd1 _3269_/A sky130_fd_sc_hd__clkbuf_4
X_3203_ _3695_/Q _3201_/Y _3202_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2401__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3134_ _3826_/Q _3134_/B _3134_/C vssd1 vssd1 vccd1 vccd1 _3134_/Y sky130_fd_sc_hd__nand3_1
X_3065_ _3123_/A _3065_/B vssd1 vssd1 vccd1 vccd1 _3065_/Y sky130_fd_sc_hd__nand2b_1
X_2016_ _3765_/Q _3749_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _4111_/CLK _3967_/D vssd1 vssd1 vccd1 vccd1 _3967_/Q sky130_fd_sc_hd__dfxtp_1
X_2918_ _2937_/A _2918_/B _2918_/C _2918_/D vssd1 vssd1 vccd1 vccd1 _2919_/B sky130_fd_sc_hd__or4_1
XANTENNA__2242__C1 _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3898_ _3902_/CLK _3898_/D vssd1 vssd1 vccd1 vccd1 _3898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2849_ _3656_/A _2849_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__and3_1
Xhold130 _3683_/X vssd1 vssd1 vccd1 vccd1 _4113_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _3981_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _3606_/X vssd1 vssd1 vccd1 vccd1 _4051_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _3406_/X vssd1 vssd1 vccd1 vccd1 _3968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _3961_/Q vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _3947_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _3446_/X vssd1 vssd1 vccd1 vccd1 _4001_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2848__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout66_A _2232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output47_A _3813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3264__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2075__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3821_ _3860_/CLK _3821_/D vssd1 vssd1 vccd1 vccd1 _3821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3752_ _3767_/CLK _3752_/D vssd1 vssd1 vccd1 vccd1 _3752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _1868_/Y hold129/X _3683_/S vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2703_ _2671_/X _2690_/Y _2702_/X vssd1 vssd1 vccd1 vccd1 _3726_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2634_ _2637_/B _2637_/C vssd1 vssd1 vccd1 vccd1 _2634_/Y sky130_fd_sc_hd__xnor2_1
X_2565_ _3720_/Q _2562_/Y _2564_/Y _2558_/Y _2560_/Y vssd1 vssd1 vccd1 vccd1 _2565_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__1943__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2496_ hold43/A _3996_/Q _4012_/Q hold61/A _2582_/S1 _2582_/S0 vssd1 vssd1 vccd1
+ vccd1 _2496_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3117_ _3199_/A hold699/X _3199_/B vssd1 vssd1 vccd1 vccd1 _3117_/X sky130_fd_sc_hd__a21o_1
X_4097_ _4105_/CLK _4097_/D vssd1 vssd1 vccd1 vccd1 _4097_/Q sky130_fd_sc_hd__dfxtp_1
X_3048_ _3048_/A _3048_/B vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3544__S _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout80 _1862_/Y vssd1 vssd1 vccd1 vccd1 _3633_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout91 _3467_/A vssd1 vssd1 vccd1 vccd1 _3320_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3902_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2350_ _2350_/A _2350_/B vssd1 vssd1 vccd1 vccd1 _2352_/B sky130_fd_sc_hd__or2_1
X_2281_ _4083_/Q _2281_/B vssd1 vssd1 vccd1 vccd1 _2338_/B sky130_fd_sc_hd__xnor2_2
X_4020_ _4029_/CLK _4020_/D vssd1 vssd1 vccd1 vccd1 _4020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1996_ hold300/X hold265/X _1996_/S vssd1 vssd1 vccd1 vccd1 _2327_/B sky130_fd_sc_hd__mux2_4
X_3804_ _4095_/CLK _3804_/D vssd1 vssd1 vccd1 vccd1 _3804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3735_ _3803_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
X_3666_ _2378_/A hold589/X _3674_/S vssd1 vssd1 vccd1 vccd1 _4097_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2617_ _2733_/S _2734_/S vssd1 vssd1 vccd1 vccd1 _3589_/A sky130_fd_sc_hd__nand2b_4
X_3597_ _4046_/Q _3592_/B _2621_/A vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2548_ hold688/X _2535_/X _2547_/X _2534_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3693_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2479_ _2612_/B _2463_/X _2465_/X _2478_/X vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3219__A1 _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1850_ _4017_/Q vssd1 vssd1 vccd1 vccd1 _3472_/A sky130_fd_sc_hd__inv_2
XFILLER_0_71_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3520_ _3520_/A _3520_/B vssd1 vssd1 vccd1 vccd1 _3520_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 _3919_/Q vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _3920_/Q vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1953__A1 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3451_ _3637_/A0 hold203/X _3453_/S vssd1 vssd1 vccd1 vccd1 _3451_/X sky130_fd_sc_hd__mux2_1
Xhold729 _4026_/Q vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_3382_ _3637_/A0 hold157/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3382_/X sky130_fd_sc_hd__mux2_1
X_2402_ _2564_/A _2402_/B vssd1 vssd1 vccd1 vccd1 _2402_/Y sky130_fd_sc_hd__nand2b_1
X_2333_ _2349_/B _2332_/X _3540_/A vssd1 vssd1 vccd1 vccd1 _2333_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2264_ _2208_/B _2148_/X _2194_/A vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4003_ _4011_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2195_ _2222_/A _2221_/B _2221_/C _2194_/Y _2220_/B vssd1 vssd1 vccd1 vccd1 _2195_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3091__C1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3394__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1979_ _1979_/A _1996_/S vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3718_ _4072_/CLK _3718_/D vssd1 vssd1 vccd1 vccd1 _3718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3649_ _2664_/X _3640_/X _3648_/X vssd1 vssd1 vccd1 vccd1 _4085_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2672__A2 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 hold615/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2951_ hold544/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2951_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2591__B _2592_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4029_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1902_ _3602_/A _3600_/B _1902_/C vssd1 vssd1 vccd1 vccd1 _1902_/X sky130_fd_sc_hd__or3_2
X_2882_ _2667_/X _2871_/X _2881_/X vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold515 _3743_/Q vssd1 vssd1 vccd1 vccd1 _2750_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _3507_/A _2277_/B _3502_/X vssd1 vssd1 vccd1 vccd1 _3505_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold526 _2764_/X vssd1 vssd1 vccd1 vccd1 _3748_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold504 _3784_/Q vssd1 vssd1 vccd1 vccd1 _2845_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _2950_/Y vssd1 vssd1 vccd1 vccd1 _3813_/D sky130_fd_sc_hd__buf_1
Xhold537 _2948_/Y vssd1 vssd1 vccd1 vccd1 _3812_/D sky130_fd_sc_hd__clkdlybuf4s25_1
X_3434_ _3682_/A0 hold67/X _3435_/S vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__mux2_1
Xhold559 _3695_/Q vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__clkbuf_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _2661_/X _3358_/X _3364_/X vssd1 vssd1 vccd1 vccd1 _3939_/D sky130_fd_sc_hd__a21o_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2362_/S _3558_/B vssd1 vssd1 vccd1 vccd1 _2316_/X sky130_fd_sc_hd__or2_1
X_3296_ _3601_/A _3296_/B vssd1 vssd1 vccd1 vccd1 _3914_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2356_/B _4085_/Q vssd1 vssd1 vccd1 vccd1 _2247_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2178_ _2178_/A _2178_/B vssd1 vssd1 vccd1 vccd1 _2179_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2590__A1 hold559/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput24 _1976_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput46 _3812_/Q vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_12
XANTENNA_fanout96_A _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput35 _1889_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3150_ _3157_/A _3150_/B vssd1 vssd1 vccd1 vccd1 _3150_/Y sky130_fd_sc_hd__nor2_1
X_3081_ _3081_/A _3090_/C vssd1 vssd1 vccd1 vccd1 _3081_/Y sky130_fd_sc_hd__nor2_1
X_2101_ _2097_/X _2100_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2101_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2078__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2032_ _3739_/Q _3796_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2032_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3983_ _4016_/CLK _3983_/D vssd1 vssd1 vccd1 vccd1 _3983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2934_ _3829_/Q _3099_/C _3100_/A vssd1 vssd1 vccd1 vccd1 _3132_/A sky130_fd_sc_hd__or3b_1
X_2865_ _2869_/A _2865_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__and3_1
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold301 _2929_/X vssd1 vssd1 vccd1 vccd1 _3805_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2796_ _2678_/X _2779_/X _2795_/X vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__a21o_1
Xhold334 hold745/X vssd1 vssd1 vccd1 vccd1 _1846_/A sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold323 _3064_/Y vssd1 vssd1 vccd1 vccd1 _3831_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _4093_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _3823_/Q vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__clkbuf_2
Xhold367 _4048_/Q vssd1 vssd1 vccd1 vccd1 _2009_/A sky130_fd_sc_hd__clkbuf_2
Xhold345 _3870_/Q vssd1 vssd1 vccd1 vccd1 _2408_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _3944_/Q vssd1 vssd1 vccd1 vccd1 _3374_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ _3675_/A _3445_/A vssd1 vssd1 vccd1 vccd1 _3425_/S sky130_fd_sc_hd__or2_4
Xhold389 _3759_/Q vssd1 vssd1 vccd1 vccd1 _2787_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2777__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3348_ _3352_/A _3348_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3348_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ input5/X hold634/X _3283_/S vssd1 vssd1 vccd1 vccd1 _3279_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2650_ _2296_/B _2737_/B _2677_/B vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__a21o_1
X_2581_ _2585_/A _2580_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3202_ _1889_/Y _3201_/A _2410_/B _2407_/D vssd1 vssd1 vccd1 vccd1 _3202_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2401__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3133_ _3133_/A _3133_/B vssd1 vssd1 vccd1 vccd1 _3136_/B sky130_fd_sc_hd__nor2_1
X_3064_ _2923_/B _2922_/Y _3063_/Y vssd1 vssd1 vccd1 vccd1 _3064_/Y sky130_fd_sc_hd__a21oi_1
X_2015_ _2013_/X _2014_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3966_ _4111_/CLK _3966_/D vssd1 vssd1 vccd1 vccd1 _3966_/Q sky130_fd_sc_hd__dfxtp_1
X_2917_ _3571_/A _3488_/A _3881_/Q _1845_/Y _2907_/X vssd1 vssd1 vccd1 vccd1 _2918_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ _4080_/CLK _3897_/D vssd1 vssd1 vccd1 vccd1 _3897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2848_ _2671_/X _2835_/Y _2847_/X vssd1 vssd1 vccd1 vccd1 _3785_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2779_ _3322_/A _2872_/A vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__and2_2
Xhold131 _3960_/Q vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _3422_/X vssd1 vssd1 vccd1 vccd1 _3981_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _3255_/X vssd1 vssd1 vccd1 vccd1 _3896_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _3974_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _3399_/X vssd1 vssd1 vccd1 vccd1 _3961_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _4074_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _3379_/X vssd1 vssd1 vccd1 vccd1 _3947_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _3966_/Q vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2784__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3860_/CLK _3820_/D vssd1 vssd1 vccd1 vccd1 _3820_/Q sky130_fd_sc_hd__dfxtp_1
X_3751_ _3767_/CLK _3751_/D vssd1 vssd1 vccd1 vccd1 _3751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2702_ _3656_/A _2702_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2702_/X sky130_fd_sc_hd__and3_1
X_3682_ _3682_/A0 hold21/X _3683_/S vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
XFILLER_0_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2633_ _2630_/A _2640_/B _2632_/Y _3227_/A vssd1 vssd1 vccd1 vccd1 _3705_/D sky130_fd_sc_hd__o211a_1
X_2564_ _2564_/A _2564_/B vssd1 vssd1 vccd1 vccd1 _2564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1943__B _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2495_ _2564_/A _2495_/B vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3116_ _2937_/A _3307_/B _3275_/C vssd1 vssd1 vccd1 vccd1 _3116_/X sky130_fd_sc_hd__a21o_1
X_4096_ _4101_/CLK _4096_/D vssd1 vssd1 vccd1 vccd1 _4096_/Q sky130_fd_sc_hd__dfxtp_1
X_3047_ _4020_/Q _3047_/B vssd1 vssd1 vccd1 vccd1 _3053_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2463__B1 _3551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2766__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3949_ _4081_/CLK _3949_/D vssd1 vssd1 vccd1 vccd1 _3949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2176__S _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout81 _1861_/Y vssd1 vssd1 vccd1 vccd1 _3676_/A0 sky130_fd_sc_hd__buf_4
Xfanout92 _3467_/A vssd1 vssd1 vccd1 vccd1 _3247_/A sky130_fd_sc_hd__buf_2
XANTENNA__2757__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout70 _2153_/S vssd1 vssd1 vccd1 vccd1 _2157_/S sky130_fd_sc_hd__buf_4
XFILLER_0_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2280_ _4082_/Q _2280_/B vssd1 vssd1 vccd1 vccd1 _2345_/S sky130_fd_sc_hd__and2_1
XANTENNA__2875__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2540__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1938__B _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ _3803_/CLK _3803_/D vssd1 vssd1 vccd1 vccd1 _3803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1995_ _2194_/A vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3734_ _3803_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_3665_ _2421_/A hold330/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__mux2_1
X_2616_ _2616_/A _2616_/B _2616_/C vssd1 vssd1 vccd1 vccd1 _2734_/S sky130_fd_sc_hd__or3_4
X_3596_ _3596_/A _3596_/B vssd1 vssd1 vccd1 vccd1 _3596_/Y sky130_fd_sc_hd__nor2_1
X_2547_ _2393_/B _2546_/X _2535_/X vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__a21bo_1
X_2478_ _2393_/B _2477_/X _2466_/X vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__a21bo_1
X_4079_ _4080_/CLK _4079_/D vssd1 vssd1 vccd1 vccd1 _4079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1864__A _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold719 _3319_/X vssd1 vssd1 vccd1 vccd1 _3320_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold708 _3314_/X vssd1 vssd1 vccd1 vccd1 _3315_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3450_ _3636_/A0 hold109/X _3453_/S vssd1 vssd1 vccd1 vccd1 _3450_/X sky130_fd_sc_hd__mux2_1
X_2401_ _3977_/Q hold55/A _3961_/Q hold75/A _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2402_/B sky130_fd_sc_hd__mux4_1
X_3381_ _3636_/A0 hold243/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3381_/X sky130_fd_sc_hd__mux2_1
X_2332_ _2306_/A _2234_/B _2331_/X vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4002_ _4011_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
X_2263_ _2031_/X _2208_/C _1995_/Y vssd1 vssd1 vccd1 vccd1 _2263_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2194_ _2194_/A _2194_/B vssd1 vssd1 vccd1 vccd1 _2194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1978_ _2230_/A _1978_/B vssd1 vssd1 vccd1 vccd1 _2392_/A sky130_fd_sc_hd__nand2_4
X_3717_ _4072_/CLK _3717_/D vssd1 vssd1 vccd1 vccd1 _3717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3648_ _3654_/A _3648_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3579_ _4042_/Q _3579_/B vssd1 vssd1 vccd1 vccd1 _3579_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4105_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2950_ _3635_/A0 _2940_/X _2949_/Y vssd1 vssd1 vccd1 vccd1 _2950_/Y sky130_fd_sc_hd__a21oi_1
X_2881_ _2887_/A _2881_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2881_/X sky130_fd_sc_hd__and3_1
X_1901_ _1895_/A _1895_/B _1899_/A _1899_/B vssd1 vssd1 vccd1 vccd1 _1987_/A sky130_fd_sc_hd__a211o_2
XFILLER_0_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3502_ _3506_/A _3502_/B vssd1 vssd1 vccd1 vccd1 _3502_/X sky130_fd_sc_hd__xor2_2
Xhold527 _3771_/Q vssd1 vssd1 vccd1 vccd1 _2813_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _3901_/Q vssd1 vssd1 vccd1 vccd1 _3265_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold505 _2846_/X vssd1 vssd1 vccd1 vccd1 _3784_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _3637_/A0 hold215/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3433_/X sky130_fd_sc_hd__mux2_1
Xhold549 _3857_/Q vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _3928_/Q vssd1 vssd1 vccd1 vccd1 _3338_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3656_/A _3364_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3364_/X sky130_fd_sc_hd__and3_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ input4/X hold651/X _3301_/S vssd1 vssd1 vccd1 vccd1 _3296_/B sky130_fd_sc_hd__mux2_1
X_2315_ _3554_/A _2315_/B vssd1 vssd1 vccd1 vccd1 _3558_/B sky130_fd_sc_hd__nor2_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2285_/B vssd1 vssd1 vccd1 vccd1 _2246_/Y sky130_fd_sc_hd__inv_2
X_2177_ _2178_/A _2178_/B vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3367__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput25 _4122_/X vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput47 _3813_/Q vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput36 _3837_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
XANTENNA_fanout89_A _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3080_ _3088_/A _3080_/B vssd1 vssd1 vccd1 vccd1 _3090_/C sky130_fd_sc_hd__nand2_1
X_2100_ _2098_/X _2099_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2100_/X sky130_fd_sc_hd__mux2_1
X_2031_ _2194_/B _2192_/B _2192_/C vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__or3_1
XANTENNA__2883__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3982_ _4111_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ _1979_/A _2925_/Y _2932_/X _3601_/A vssd1 vssd1 vccd1 vccd1 _2933_/X sky130_fd_sc_hd__o211a_1
X_2864_ _2667_/X _2853_/X _2863_/X vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3349__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2795_ _2813_/A _2795_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2795_/X sky130_fd_sc_hd__and3_1
Xhold302 _3847_/Q vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold324 hold735/X vssd1 vssd1 vccd1 vccd1 _2642_/A sky130_fd_sc_hd__buf_1
Xhold335 _3228_/X vssd1 vssd1 vccd1 vccd1 _3229_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _3662_/X vssd1 vssd1 vccd1 vccd1 _4093_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _2995_/Y vssd1 vssd1 vccd1 vccd1 _3823_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _2646_/D vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__clkbuf_4
Xhold346 _3217_/X vssd1 vssd1 vccd1 vccd1 _3870_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _3846_/Q vssd1 vssd1 vccd1 vccd1 _3165_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3416_ _3639_/A0 hold211/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3416_/X sky130_fd_sc_hd__mux2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ _2661_/X _3340_/X _3346_/X vssd1 vssd1 vccd1 vccd1 _3931_/D sky130_fd_sc_hd__a21o_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3601_/A _3278_/B vssd1 vssd1 vccd1 vccd1 _3906_/D sky130_fd_sc_hd__and2_1
XANTENNA__2088__A1 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2229_ _2424_/B _2229_/B vssd1 vssd1 vccd1 vccd1 _2230_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2580_ hold69/A hold77/A _4016_/Q hold81/A _2584_/S1 _2582_/S0 vssd1 vssd1 vccd1
+ vccd1 _2580_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3503__A1 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2089__S _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3201_ _3201_/A _3201_/B vssd1 vssd1 vccd1 vccd1 _3201_/Y sky130_fd_sc_hd__nand2_2
X_3132_ _3132_/A _3132_/B vssd1 vssd1 vccd1 vccd1 _3133_/B sky130_fd_sc_hd__nor2_1
X_3063_ _2923_/B _2922_/Y _3601_/A vssd1 vssd1 vccd1 vccd1 _3063_/Y sky130_fd_sc_hd__o21ai_1
X_2014_ _3741_/Q _3757_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3502__A _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _4113_/CLK _3965_/D vssd1 vssd1 vccd1 vccd1 _3965_/Q sky130_fd_sc_hd__dfxtp_1
X_2916_ _4035_/Q _1856_/Y _1860_/Y _4031_/Q _2915_/X vssd1 vssd1 vccd1 vccd1 _2918_/C
+ sky130_fd_sc_hd__a221o_1
X_3896_ _4072_/CLK _3896_/D vssd1 vssd1 vccd1 vccd1 _3896_/Q sky130_fd_sc_hd__dfxtp_1
X_2847_ _3269_/A _2847_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2847_/X sky130_fd_sc_hd__and3_1
Xhold110 _3450_/X vssd1 vssd1 vccd1 vccd1 _4005_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2778_ _2678_/X _2761_/X _2777_/X vssd1 vssd1 vccd1 vccd1 _2778_/X sky130_fd_sc_hd__a21o_1
Xhold132 _3396_/X vssd1 vssd1 vccd1 vccd1 _3960_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _3994_/Q vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _3967_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _3632_/X vssd1 vssd1 vccd1 vccd1 _4074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _3414_/X vssd1 vssd1 vccd1 vccd1 _3974_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _3969_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _3404_/X vssd1 vssd1 vccd1 vccd1 _3966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _4067_/Q vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3430__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2698__A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3249__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3322__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3421__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3750_ _3791_/CLK _3750_/D vssd1 vssd1 vccd1 vccd1 _3750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2701_ _2667_/X _2690_/Y _2700_/X vssd1 vssd1 vccd1 vccd1 _3725_/D sky130_fd_sc_hd__a21o_1
X_3681_ _1866_/Y hold171/X _3683_/S vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2632_ _2640_/B _2632_/B vssd1 vssd1 vccd1 vccd1 _2632_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2563_ hold83/A _3896_/Q _3702_/Q hold89/A _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2564_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2494_ hold65/A _4069_/Q _4061_/Q hold71/A _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2495_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3115_ _3133_/A _3115_/B vssd1 vssd1 vccd1 vccd1 _3307_/B sky130_fd_sc_hd__nand2b_1
X_4095_ _4095_/CLK _4095_/D vssd1 vssd1 vccd1 vccd1 _4095_/Q sky130_fd_sc_hd__dfxtp_1
X_3046_ _4018_/Q _3046_/B vssd1 vssd1 vccd1 vccd1 _3052_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__2999__C1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2463__A1 _2232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3660__A0 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3412__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3948_ _4080_/CLK _3948_/D vssd1 vssd1 vccd1 vccd1 _3948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3879_ _4031_/CLK _3879_/D vssd1 vssd1 vccd1 vccd1 _3879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3403__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout60 _2155_/S vssd1 vssd1 vccd1 vccd1 _2119_/S sky130_fd_sc_hd__buf_6
Xfanout82 hold663/X vssd1 vssd1 vccd1 vccd1 _3602_/A sky130_fd_sc_hd__clkbuf_8
Xfanout71 _1919_/Y vssd1 vssd1 vccd1 vccd1 _2153_/S sky130_fd_sc_hd__buf_4
Xfanout93 _3114_/A vssd1 vssd1 vccd1 vccd1 _3131_/A sky130_fd_sc_hd__buf_4
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4042_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output52_A _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2693__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2540__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ _4047_/CLK _3802_/D vssd1 vssd1 vccd1 vccd1 _3802_/Q sky130_fd_sc_hd__dfxtp_1
X_1994_ _2142_/A _3554_/B _1993_/X _1988_/A vssd1 vssd1 vccd1 vccd1 _2194_/A sky130_fd_sc_hd__o22a_4
XFILLER_0_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3733_ _4047_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3664_ _2327_/B hold265/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2615_ _2733_/S _2615_/B vssd1 vssd1 vccd1 vccd1 _2640_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3595_ _3592_/A _2613_/Y _3593_/X _3594_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _4046_/D
+ sky130_fd_sc_hd__o221a_1
X_2546_ _2545_/X input10/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__mux2_1
X_2477_ _2476_/X input13/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__mux2_1
X_4078_ _4081_/CLK _4078_/D vssd1 vssd1 vccd1 vccd1 _4078_/Q sky130_fd_sc_hd__dfxtp_1
X_3029_ _3856_/Q _3032_/A vssd1 vssd1 vccd1 vccd1 _3030_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3633__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3624__A0 _1862_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold709 _3832_/Q vssd1 vssd1 vccd1 vccd1 _3123_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2400_ _2564_/A _2399_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2400_/Y sky130_fd_sc_hd__a21oi_1
X_3380_ _3635_/A0 hold227/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3380_/X sky130_fd_sc_hd__mux2_1
X_2331_ _2737_/C _2285_/X _2329_/X _2330_/X vssd1 vssd1 vccd1 vccd1 _2331_/X sky130_fd_sc_hd__a31o_1
X_2262_ _2005_/B _2220_/B _2093_/B _2207_/X vssd1 vssd1 vccd1 vccd1 _2266_/B sky130_fd_sc_hd__a211oi_2
XANTENNA__2097__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _4014_/CLK _4001_/D vssd1 vssd1 vccd1 vccd1 _4001_/Q sky130_fd_sc_hd__dfxtp_1
X_2193_ _3693_/Q _2048_/S _2084_/X _2194_/B vssd1 vssd1 vccd1 vccd1 _2221_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3615__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3716_ _3905_/CLK _3716_/D vssd1 vssd1 vccd1 vccd1 _3716_/Q sky130_fd_sc_hd__dfxtp_1
X_1977_ _2646_/B _1977_/B vssd1 vssd1 vccd1 vccd1 _2512_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3647_ _2661_/X _3640_/X _3646_/X vssd1 vssd1 vccd1 vccd1 _4084_/D sky130_fd_sc_hd__a21o_1
X_3578_ hold1/X _2646_/D _3577_/X _3587_/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o211a_1
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2529_ _2431_/Y _2529_/B _2571_/C vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__and3b_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3606__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2440__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2880_ _2664_/X _2871_/X _2879_/X vssd1 vssd1 vccd1 vccd1 _3799_/D sky130_fd_sc_hd__a21o_1
XANTENNA__2820__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1900_ _1895_/A _1895_/B _1899_/A _1899_/B vssd1 vssd1 vccd1 vccd1 _1906_/A sky130_fd_sc_hd__a211oi_4
XFILLER_0_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3501_ hold581/X _3564_/B _3499_/Y _3500_/X _3587_/A vssd1 vssd1 vccd1 vccd1 _3501_/X
+ sky130_fd_sc_hd__o221a_1
Xhold517 _3793_/Q vssd1 vssd1 vccd1 vccd1 _2865_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 _3922_/Q vssd1 vssd1 vccd1 vccd1 _3326_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _3636_/A0 hold53/X _3435_/S vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__mux2_1
Xhold528 _2814_/X vssd1 vssd1 vccd1 vccd1 _3771_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _3339_/X vssd1 vssd1 vccd1 vccd1 _3928_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _2658_/X _3358_/X _3362_/X vssd1 vssd1 vccd1 vccd1 _3938_/D sky130_fd_sc_hd__a21o_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2313_/A _2313_/B _2349_/B vssd1 vssd1 vccd1 vccd1 _2314_/X sky130_fd_sc_hd__a21o_1
X_3294_ _3294_/A _3294_/B vssd1 vssd1 vccd1 vccd1 _3301_/S sky130_fd_sc_hd__nand2_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _4085_/Q _2356_/B vssd1 vssd1 vccd1 vccd1 _2285_/B sky130_fd_sc_hd__and2b_1
X_2176_ _2606_/A _2175_/Y _3544_/S vssd1 vssd1 vccd1 vccd1 _2178_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2498__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput48 _3814_/Q vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__buf_12
Xoutput26 _1973_/X vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__buf_12
Xoutput37 _3918_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
XANTENNA__2878__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2802__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2030_ _2256_/A _2165_/B _3502_/B vssd1 vssd1 vccd1 vccd1 _2192_/C sky130_fd_sc_hd__and3_1
X_3981_ _4113_/CLK _3981_/D vssd1 vssd1 vccd1 vccd1 _3981_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2932_ input7/X _3834_/Q _3072_/B vssd1 vssd1 vccd1 vccd1 _2932_/X sky130_fd_sc_hd__or3_1
X_2863_ _2863_/A _2863_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2794_ _2674_/X _2779_/X _2793_/X vssd1 vssd1 vccd1 vccd1 _3762_/D sky130_fd_sc_hd__a21o_1
Xhold325 _3580_/X vssd1 vssd1 vccd1 vccd1 _4042_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold303 _3168_/X vssd1 vssd1 vccd1 vccd1 _3847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _3869_/Q vssd1 vssd1 vccd1 vccd1 _2408_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _4014_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _4009_/Q vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _3572_/X vssd1 vssd1 vccd1 vccd1 _4038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _3868_/Q vssd1 vssd1 vccd1 vccd1 _2408_/C sky130_fd_sc_hd__dlygate4sd3_1
X_3415_ _3682_/A0 hold223/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3415_/X sky130_fd_sc_hd__mux2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _3656_/A _3346_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3346_/X sky130_fd_sc_hd__and3_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ input4/X hold683/X _3283_/S vssd1 vssd1 vccd1 vccd1 _3278_/B sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _2378_/A _2378_/B vssd1 vssd1 vccd1 vccd1 _2229_/B sky130_fd_sc_hd__and2_1
X_2159_ _3715_/Q _3727_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2160_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3200_ _2957_/Y _3199_/X _3114_/A vssd1 vssd1 vccd1 vccd1 _3862_/D sky130_fd_sc_hd__o21a_1
X_3131_ _3131_/A _3131_/B vssd1 vssd1 vccd1 vccd1 _3837_/D sky130_fd_sc_hd__and2_1
X_3062_ _3320_/A _3062_/B vssd1 vssd1 vccd1 vccd1 _3830_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2013_ hold47/A _3797_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ _4111_/CLK _3964_/D vssd1 vssd1 vccd1 vccd1 _3964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2915_ _1841_/Y _3885_/Q _3883_/Q _1843_/Y vssd1 vssd1 vccd1 vccd1 _2915_/X sky130_fd_sc_hd__a22o_1
X_3895_ _4081_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2846_ _2667_/X _2835_/Y _2845_/X vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__a21o_1
X_2777_ _2813_/A _2777_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2777_/X sky130_fd_sc_hd__and3_1
Xhold100 _3384_/X vssd1 vssd1 vccd1 vccd1 _3952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _3438_/X vssd1 vssd1 vccd1 vccd1 _3994_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _3405_/X vssd1 vssd1 vccd1 vccd1 _3967_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _3958_/Q vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold133 _3897_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _4070_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _3892_/Q vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _3409_/X vssd1 vssd1 vccd1 vccd1 _3969_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold199 _4075_/Q vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _3624_/X vssd1 vssd1 vccd1 vccd1 _4067_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _2661_/X _3322_/X _3328_/X vssd1 vssd1 vccd1 vccd1 _3923_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1992__A1 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2979__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2941__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2700_ _3269_/A _2700_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__and3_1
X_3680_ _1865_/Y hold251/X _3683_/S vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xload_slew1 _1906_/A vssd1 vssd1 vccd1 vccd1 _1988_/A sky130_fd_sc_hd__buf_2
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _3589_/A _2637_/C _2630_/Y _2734_/S _2142_/A vssd1 vssd1 vccd1 vccd1 _2631_/X
+ sky130_fd_sc_hd__o32a_1
X_2562_ _3719_/Q _2562_/B vssd1 vssd1 vccd1 vccd1 _2562_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2493_ _2392_/X _2485_/X _2391_/X vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3513__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3114_ _3114_/A _3114_/B vssd1 vssd1 vccd1 vccd1 _3836_/D sky130_fd_sc_hd__and2_1
X_4094_ _4101_/CLK _4094_/D vssd1 vssd1 vccd1 vccd1 _4094_/Q sky130_fd_sc_hd__dfxtp_1
X_3045_ _3850_/Q _3849_/Q vssd1 vssd1 vccd1 vccd1 _3046_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3947_ _4095_/CLK _3947_/D vssd1 vssd1 vccd1 vccd1 _3947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3878_ _4014_/CLK _3878_/D vssd1 vssd1 vccd1 vccd1 _3878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2829_ _2869_/A _2829_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__and3_1
XANTENNA__2799__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout72 _2151_/S vssd1 vssd1 vccd1 vccd1 _2158_/S sky130_fd_sc_hd__clkbuf_8
Xfanout61 _1930_/Y vssd1 vssd1 vccd1 vccd1 _3544_/S sky130_fd_sc_hd__buf_4
Xfanout83 hold663/X vssd1 vssd1 vccd1 vccd1 _2008_/C sky130_fd_sc_hd__buf_2
Xfanout94 _3658_/B vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3801_ _4047_/CLK _3801_/D vssd1 vssd1 vccd1 vccd1 _3801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1993_ _2151_/S _1992_/X _3544_/S vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3732_ _4045_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3663_ _3540_/A hold636/X _3674_/S vssd1 vssd1 vccd1 vccd1 _4094_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2614_ _2614_/A _2614_/B vssd1 vssd1 vccd1 vccd1 _2615_/B sky130_fd_sc_hd__or2_2
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3594_ _3529_/A _3589_/A _2615_/B vssd1 vssd1 vccd1 vccd1 _3594_/X sky130_fd_sc_hd__a21o_1
X_2545_ _1882_/Y _2544_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2545_/X sky130_fd_sc_hd__mux2_1
X_2476_ _1885_/Y _2475_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__mux2_1
X_4077_ _4077_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
X_3028_ _4025_/Q _3028_/B vssd1 vssd1 vccd1 vccd1 _3056_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2675__A2 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2330_ _1945_/Y _2233_/X _2235_/Y _2616_/A _2181_/Y vssd1 vssd1 vccd1 vccd1 _2330_/X
+ sky130_fd_sc_hd__o221a_1
X_2261_ _4084_/Q _2604_/B _2261_/C vssd1 vssd1 vccd1 vccd1 _2350_/B sky130_fd_sc_hd__and3_1
X_4000_ _4016_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2192_ _2192_/A _2192_/B _2192_/C vssd1 vssd1 vccd1 vccd1 _2221_/B sky130_fd_sc_hd__or3_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3379__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ _3602_/A _1978_/B vssd1 vssd1 vccd1 vccd1 _1976_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3715_ _3795_/CLK _3715_/D vssd1 vssd1 vccd1 vccd1 _3715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2142__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _3656_/A _3646_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__and3_1
X_3577_ _4041_/Q _3579_/B vssd1 vssd1 vccd1 vccd1 _3577_/X sky130_fd_sc_hd__or2_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2354__A1 _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2528_ _2570_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2529_/B sky130_fd_sc_hd__nor2_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _2571_/B _2550_/B _2571_/C vssd1 vssd1 vccd1 vccd1 _2459_/X sky130_fd_sc_hd__a21o_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2345__A1 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2440__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2661__S _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _3584_/A _3554_/B hold368/X vssd1 vssd1 vccd1 vccd1 _3500_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold518 hold741/X vssd1 vssd1 vccd1 vccd1 _1843_/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold507 _3713_/Q vssd1 vssd1 vccd1 vccd1 _2666_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3431_ _3635_/A0 hold61/X _3435_/S vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__mux2_1
Xhold529 _3789_/Q vssd1 vssd1 vccd1 vccd1 _2857_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3654_/A _3362_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3362_/X sky130_fd_sc_hd__and3_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2313_/A _2313_/B vssd1 vssd1 vccd1 vccd1 _2435_/A sky130_fd_sc_hd__and2_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3658_/B _3293_/B vssd1 vssd1 vccd1 vccd1 _3913_/D sky130_fd_sc_hd__and2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2232_/S _3529_/B _2242_/X vssd1 vssd1 vccd1 vccd1 _2356_/B sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4011_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2175_ _2175_/A vssd1 vssd1 vccd1 vccd1 _2175_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2498__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1959_ _2230_/A _2158_/S _1959_/C _1959_/D vssd1 vssd1 vccd1 vccd1 _2647_/A sky130_fd_sc_hd__and4_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3629_ _3682_/A0 hold167/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3629_/X sky130_fd_sc_hd__mux2_1
Xoutput49 _3815_/Q vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__buf_12
Xoutput27 _4123_/X vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__buf_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput38 _3919_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
XFILLER_0_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3980_ _4111_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _1989_/A _2925_/Y _2930_/X _3601_/A vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2862_ _2664_/X _2853_/X _2861_/X vssd1 vssd1 vccd1 vccd1 _3791_/D sky130_fd_sc_hd__a21o_1
X_2793_ _2805_/A _2793_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__and3_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold326 _3838_/Q vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _3804_/Q vssd1 vssd1 vccd1 vccd1 _1925_/C sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold315 _3215_/X vssd1 vssd1 vccd1 vccd1 _3869_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2309__A1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold348 _3466_/X vssd1 vssd1 vccd1 vccd1 _3467_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2309__B2 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3414_ _3637_/A0 hold153/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3414_/X sky130_fd_sc_hd__mux2_1
Xhold337 _3213_/X vssd1 vssd1 vccd1 vccd1 _3868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 _3456_/X vssd1 vssd1 vccd1 vccd1 _3457_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _2658_/X _3340_/X _3344_/X vssd1 vssd1 vccd1 vccd1 _3930_/D sky130_fd_sc_hd__a21o_1
X_3276_ _3276_/A _3276_/B _3285_/D vssd1 vssd1 vccd1 vccd1 _3283_/S sky130_fd_sc_hd__or3_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2226_/X _3540_/B _2227_/S vssd1 vssd1 vccd1 vccd1 _2227_/X sky130_fd_sc_hd__mux2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _2156_/X _2157_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2158_/X sky130_fd_sc_hd__mux2_1
X_2089_ _2119_/S _2088_/X _3544_/S vssd1 vssd1 vccd1 vccd1 _2089_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2796__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout94_A _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3130_ hold712/X _3129_/X _3130_/S vssd1 vssd1 vccd1 vccd1 _3130_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3071__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3061_ _3100_/A _3065_/B _3008_/X _3060_/Y vssd1 vssd1 vccd1 vccd1 _3062_/B sky130_fd_sc_hd__o2bb2a_1
X_2012_ _2256_/A _2165_/B vssd1 vssd1 vccd1 vccd1 _2048_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3963_ _4112_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2778__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2914_ _4041_/Q _1853_/Y _3884_/Q _1842_/Y _2913_/X vssd1 vssd1 vccd1 vccd1 _2919_/A
+ sky130_fd_sc_hd__a221o_1
X_3894_ _4081_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2845_ _3269_/A _2845_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__and3_1
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 _3957_/Q vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2776_ _2674_/X _2761_/X _2775_/X vssd1 vssd1 vccd1 vccd1 _3754_/D sky130_fd_sc_hd__a21o_1
Xhold123 _3983_/Q vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _3394_/X vssd1 vssd1 vccd1 vccd1 _3958_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _3256_/X vssd1 vssd1 vccd1 vccd1 _3897_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2950__A1 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold145 _4065_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _3627_/X vssd1 vssd1 vccd1 vccd1 _4070_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _4072_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _3698_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _3251_/X vssd1 vssd1 vccd1 vccd1 _3892_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3680__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3352_/A _3328_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__and3_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3269_/A _3259_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3259_/X sky130_fd_sc_hd__and3_1
XANTENNA__2561__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold690 _3873_/Q vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2630_ _2630_/A _2630_/B vssd1 vssd1 vccd1 vccd1 _2630_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2561_ _3983_/Q hold21/A _3967_/Q hold15/A _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2562_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2492_ _2392_/A _2489_/X _2491_/X _2612_/B vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_10_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3113_ _3112_/X hold725/X _3113_/S vssd1 vssd1 vccd1 vccd1 _3113_/X sky130_fd_sc_hd__mux2_1
X_4093_ _4101_/CLK _4093_/D vssd1 vssd1 vccd1 vccd1 _4093_/Q sky130_fd_sc_hd__dfxtp_1
X_3044_ _4019_/Q _3044_/B vssd1 vssd1 vccd1 vccd1 _3053_/A sky130_fd_sc_hd__xnor2_1
X_3946_ _4080_/CLK _3946_/D vssd1 vssd1 vccd1 vccd1 _3946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3877_ _4014_/CLK _3877_/D vssd1 vssd1 vccd1 vccd1 _3877_/Q sky130_fd_sc_hd__dfxtp_1
X_2828_ _2671_/X _2815_/X _2827_/X vssd1 vssd1 vccd1 vccd1 _3777_/D sky130_fd_sc_hd__a21o_1
X_2759_ _2678_/X _2742_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _2759_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 _1908_/X vssd1 vssd1 vccd1 vccd1 _2151_/S sky130_fd_sc_hd__clkbuf_8
Xfanout62 _2160_/A vssd1 vssd1 vccd1 vccd1 _2142_/A sky130_fd_sc_hd__clkbuf_8
Xfanout95 _3658_/B vssd1 vssd1 vccd1 vccd1 _3497_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout84 _2009_/A vssd1 vssd1 vccd1 vccd1 _3600_/B sky130_fd_sc_hd__buf_6
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2664__S _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3800_ _4042_/CLK _3800_/D vssd1 vssd1 vccd1 vccd1 _3800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3731_ _4042_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
X_1992_ _2315_/B _3506_/A _2227_/S vssd1 vssd1 vccd1 vccd1 _1992_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2602__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3862_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _3529_/A hold312/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__mux2_1
X_3593_ _3596_/B _3593_/B _3593_/C vssd1 vssd1 vccd1 vccd1 _3593_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2613_ _2614_/A _2614_/B vssd1 vssd1 vccd1 vccd1 _2613_/Y sky130_fd_sc_hd__nor2_2
X_2544_ _3720_/Q _2541_/Y _2543_/Y _2537_/Y _2539_/Y vssd1 vssd1 vccd1 vccd1 _2544_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2475_ _3720_/Q _2472_/Y _2474_/Y _2468_/Y _2470_/Y vssd1 vssd1 vccd1 vccd1 _2475_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ _4095_/CLK _4076_/D vssd1 vssd1 vccd1 vccd1 _4076_/Q sky130_fd_sc_hd__dfxtp_1
X_3027_ _3027_/A _3027_/B vssd1 vssd1 vccd1 vccd1 _3028_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3929_ _3938_/CLK _3929_/D vssd1 vssd1 vccd1 vccd1 _3929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2260_ _2604_/B _2261_/C _4084_/Q vssd1 vssd1 vccd1 vccd1 _2260_/X sky130_fd_sc_hd__a21o_1
X_2191_ _2194_/A _2191_/B _2191_/C vssd1 vssd1 vccd1 vccd1 _2191_/X sky130_fd_sc_hd__and3_1
XFILLER_0_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _3322_/A _2296_/B _3321_/A _1943_/D _1974_/B vssd1 vssd1 vccd1 vccd1 _1978_/B
+ sky130_fd_sc_hd__a41o_2
XFILLER_0_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3714_ _3905_/CLK _3714_/D vssd1 vssd1 vccd1 vccd1 _3714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3645_ _2658_/X _3640_/X _3644_/X vssd1 vssd1 vccd1 vccd1 _4083_/D sky130_fd_sc_hd__a21o_1
X_3576_ _2637_/B hold368/X hold480/X _3227_/A vssd1 vssd1 vccd1 vccd1 _4040_/D sky130_fd_sc_hd__o211a_1
XANTENNA_fanout107_A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2527_ hold609/X _2514_/Y _2526_/X _2513_/X _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3692_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2458_ _2455_/X _2457_/Y _2570_/A vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__mux2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _2392_/A _3566_/A _2382_/Y _2388_/Y vssd1 vssd1 vccd1 vccd1 _2389_/X sky130_fd_sc_hd__o31a_1
X_4059_ _4073_/CLK _4059_/D vssd1 vssd1 vccd1 vccd1 _4059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold688_A _3693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3542__A1 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2569__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold508 _2668_/X vssd1 vssd1 vccd1 vccd1 _3713_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3430_ _3634_/A0 hold79/X _3435_/S vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__mux2_1
Xhold519 _3234_/X vssd1 vssd1 vccd1 vccd1 _3235_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3361_ _2655_/X _3358_/X _3360_/X vssd1 vssd1 vccd1 vccd1 _3361_/X sky130_fd_sc_hd__a21o_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _2310_/Y _2311_/X _2309_/X vssd1 vssd1 vccd1 vccd1 _2313_/B sky130_fd_sc_hd__o21bai_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ input7/X _1949_/A _3292_/S vssd1 vssd1 vccd1 vccd1 _3292_/X sky130_fd_sc_hd__mux2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3297__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2243_ _3692_/Q _2269_/A _2200_/Y _2240_/X vssd1 vssd1 vccd1 vccd1 _3529_/B sky130_fd_sc_hd__a22o_2
X_2174_ _2170_/X _3566_/B _2227_/S vssd1 vssd1 vccd1 vccd1 _2175_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1958_ _1929_/A _1949_/X _1954_/Y _1957_/Y vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3683__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1889_ _2939_/A vssd1 vssd1 vccd1 vccd1 _1889_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3628_ _1866_/Y hold207/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3628_/X sky130_fd_sc_hd__mux2_1
Xoutput28 _4123_/A vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__buf_12
Xoutput39 _3920_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
XFILLER_0_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3559_ _3559_/A _3559_/B vssd1 vssd1 vccd1 vccd1 _3562_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3288__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3279__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3451__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2930_ input6/X _3834_/Q _3072_/B vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__or3_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2863_/A _2861_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__and3_1
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2792_ _2671_/X _2779_/X _2791_/X vssd1 vssd1 vccd1 vccd1 _3761_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold305 _2927_/X vssd1 vssd1 vccd1 vccd1 _3804_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _4090_/Q vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold327 _3139_/X vssd1 vssd1 vccd1 vccd1 _3838_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _4045_/Q vssd1 vssd1 vccd1 vccd1 _2619_/A sky130_fd_sc_hd__buf_1
Xhold338 _4103_/Q vssd1 vssd1 vccd1 vccd1 _2737_/A sky130_fd_sc_hd__buf_1
X_3413_ _3636_/A0 hold237/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3413_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1962__D _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3352_/A _3344_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3344_/X sky130_fd_sc_hd__and3_1
X_3275_ _3275_/A _3275_/B _3275_/C vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__or3_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2093_/B _2223_/X _2224_/X _2225_/X vssd1 vssd1 vccd1 vccd1 _2226_/X sky130_fd_sc_hd__a31o_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ _3935_/Q _3927_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3678__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2088_ _2268_/A _3518_/A _2227_/S vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3442__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout87_A _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3433__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2667__S _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ _3100_/A _3060_/B vssd1 vssd1 vccd1 vccd1 _3060_/Y sky130_fd_sc_hd__xnor2_1
X_2011_ _2646_/B _1978_/B _2612_/B _2737_/B vssd1 vssd1 vccd1 vccd1 _2165_/B sky130_fd_sc_hd__a31o_2
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3424__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3962_ _4113_/CLK _3962_/D vssd1 vssd1 vccd1 vccd1 _3962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2913_ _1848_/Y _4017_/Q _3880_/Q _1846_/Y _2906_/X vssd1 vssd1 vccd1 vccd1 _2913_/X
+ sky130_fd_sc_hd__a221o_1
X_3893_ _4077_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2844_ _2664_/X _2835_/Y _2843_/X vssd1 vssd1 vccd1 vccd1 _3783_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2775_ _2869_/A _2775_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__and3_1
Xhold102 _3393_/X vssd1 vssd1 vccd1 vccd1 _3957_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 _3424_/X vssd1 vssd1 vccd1 vccd1 _3983_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _3996_/Q vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _4079_/Q vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2950__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 _3621_/X vssd1 vssd1 vccd1 vccd1 _4065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _3950_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _3629_/X vssd1 vssd1 vccd1 vccd1 _4072_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _3701_/Q vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _2658_/X _3322_/X _3326_/X vssd1 vssd1 vccd1 vccd1 _3922_/D sky130_fd_sc_hd__a21o_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3258_/A _3641_/B vssd1 vssd1 vccd1 vccd1 _3273_/C sky130_fd_sc_hd__or2_2
X_3189_ _4025_/Q hold549/X _3189_/S vssd1 vssd1 vccd1 vccd1 _3189_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3663__A0 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2209_ _2222_/A _2130_/X _2148_/X _2208_/X vssd1 vssd1 vccd1 vccd1 _2209_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2561__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3415__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2941__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold680 _4044_/Q vssd1 vssd1 vccd1 vccd1 _2619_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _4087_/Q vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3406__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2560_ _2585_/A _2559_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2560_/Y sky130_fd_sc_hd__a21oi_1
X_2491_ _2512_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ hold699/X _3199_/B _3107_/X _3111_/Y vssd1 vssd1 vccd1 vccd1 _3112_/X sky130_fd_sc_hd__a2bb2o_1
X_4092_ _4092_/CLK _4092_/D vssd1 vssd1 vccd1 vccd1 _4092_/Q sky130_fd_sc_hd__dfxtp_1
X_3043_ _3043_/A _3043_/B vssd1 vssd1 vccd1 vccd1 _3044_/B sky130_fd_sc_hd__or2_1
XANTENNA__2129__C _3551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3945_ _4080_/CLK _3945_/D vssd1 vssd1 vccd1 vccd1 _3945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3876_ _4014_/CLK _3876_/D vssd1 vssd1 vccd1 vccd1 _3876_/Q sky130_fd_sc_hd__dfxtp_1
X_2827_ _2869_/A _2827_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__and3_1
X_2758_ _2813_/A _2758_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2689_ hold609/X _2681_/Y _2688_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _2689_/X sky130_fd_sc_hd__o211a_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2100__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3636__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4073_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout74 _1868_/Y vssd1 vssd1 vccd1 vccd1 _3639_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout63 _2269_/A vssd1 vssd1 vccd1 vccd1 _2230_/A sky130_fd_sc_hd__clkbuf_8
Xfanout85 _2564_/A vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__clkbuf_4
Xfanout96 _3658_/B vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3627__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2850__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3730_ _4045_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
X_1991_ hold330/X _1890_/Y _1989_/X vssd1 vssd1 vccd1 vccd1 _2421_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ _3518_/A hold257/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3661_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ _3592_/A _3592_/B vssd1 vssd1 vccd1 vccd1 _3593_/C sky130_fd_sc_hd__or2_1
X_2612_ _3658_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2614_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2543_ _2564_/A _2543_/B vssd1 vssd1 vccd1 vccd1 _2543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2474_ _2585_/A _2474_/B vssd1 vssd1 vccd1 vccd1 _2474_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3618__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3540__A _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4075_ _4080_/CLK _4075_/D vssd1 vssd1 vccd1 vccd1 _4075_/Q sky130_fd_sc_hd__dfxtp_1
X_3026_ _3856_/Q _3032_/A _3857_/Q vssd1 vssd1 vccd1 vccd1 _3027_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3928_ _3939_/CLK _3928_/D vssd1 vssd1 vccd1 vccd1 _3928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3859_ _3862_/CLK _3859_/D vssd1 vssd1 vccd1 vccd1 _3859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3609__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2832__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2596__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2190_ _3688_/Q _2048_/S _2111_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2191_/C sky130_fd_sc_hd__a211o_1
XANTENNA_output50_A _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2704__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1974_ _3201_/A _1974_/B vssd1 vssd1 vccd1 vccd1 _1977_/B sky130_fd_sc_hd__nor2_1
X_3713_ _3795_/CLK _3713_/D vssd1 vssd1 vccd1 vccd1 _3713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3644_ _3654_/A _3644_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3575_ _3575_/A _3579_/B vssd1 vssd1 vccd1 vccd1 _3575_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2526_ _2393_/B _2525_/X _2514_/Y vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__a21bo_1
X_2457_ _2549_/B vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__inv_2
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _2392_/A _2386_/X _2387_/Y _2393_/B vssd1 vssd1 vccd1 vccd1 _2388_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4058_ _4073_/CLK _4058_/D vssd1 vssd1 vccd1 vccd1 _4058_/Q sky130_fd_sc_hd__dfxtp_1
X_3009_ _3060_/B _3009_/B vssd1 vssd1 vccd1 vccd1 _3009_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2814__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 _3744_/Q vssd1 vssd1 vccd1 vccd1 _2752_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3360_ _3656_/A _3360_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3360_/X sky130_fd_sc_hd__and3_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2219_/Y _2287_/X _2308_/Y _2180_/B vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3658_/B _3291_/B vssd1 vssd1 vccd1 vccd1 _3912_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2279_/S _2240_/X _2241_/X _3544_/S vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__o211a_1
X_2173_ _2170_/X _2172_/X _3676_/A0 _2646_/B vssd1 vssd1 vccd1 vccd1 _2606_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3221__A1 _3460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1957_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1957_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1888_ _3602_/A _3600_/B vssd1 vssd1 vccd1 vccd1 _2939_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3627_ _3636_/A0 hold155/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3627_/X sky130_fd_sc_hd__mux2_1
Xoutput29 _3816_/Q vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3558_ _3558_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _3559_/B sky130_fd_sc_hd__nand2_1
X_2509_ hold609/X _2508_/C _1930_/Y vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__a21o_1
X_3489_ _3571_/A _3494_/S _3488_/Y _3587_/A vssd1 vssd1 vccd1 vccd1 _3489_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2328__B _3551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3212__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2860_ _2661_/X _2853_/X _2859_/X vssd1 vssd1 vccd1 vccd1 _3790_/D sky130_fd_sc_hd__a21o_1
XANTENNA__2254__A _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2791_ _2813_/A _2791_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__and3_1
XANTENNA__3203__A1 _3695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold306 _3807_/Q vssd1 vssd1 vccd1 vccd1 _1979_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _3659_/X vssd1 vssd1 vccd1 vccd1 _4090_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold328 _4102_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__buf_1
Xhold339 _3672_/X vssd1 vssd1 vccd1 vccd1 _4103_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _3635_/A0 hold65/X _3416_/S vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _2655_/X _3340_/X _3342_/X vssd1 vssd1 vccd1 vccd1 _3343_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _2678_/X _3257_/Y _3273_/X vssd1 vssd1 vccd1 vccd1 _3905_/D sky130_fd_sc_hd__a21o_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2094_/Y _2221_/X _2222_/X _2220_/X _2238_/B vssd1 vssd1 vccd1 vccd1 _2225_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _4088_/Q _3943_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2087_ _2221_/A _2049_/X _2086_/X vssd1 vssd1 vccd1 vccd1 _2087_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1987__B _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2989_ _3140_/C _2989_/B vssd1 vssd1 vccd1 vccd1 _2990_/C sky130_fd_sc_hd__nor2_1
XANTENNA__2953__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ _2698_/A _2616_/B _3579_/B vssd1 vssd1 vccd1 vccd1 _2737_/B sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4101_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3961_ _4111_/CLK _3961_/D vssd1 vssd1 vccd1 vccd1 _3961_/Q sky130_fd_sc_hd__dfxtp_1
X_2912_ _1839_/Y _1854_/A _3884_/Q _1842_/Y _2911_/X vssd1 vssd1 vccd1 vccd1 _2912_/X
+ sky130_fd_sc_hd__o221a_1
X_3892_ _4095_/CLK _3892_/D vssd1 vssd1 vccd1 vccd1 _3892_/Q sky130_fd_sc_hd__dfxtp_1
X_2843_ _3269_/A _2843_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__and3_1
X_2774_ _2671_/X _2761_/X _2773_/X vssd1 vssd1 vccd1 vccd1 _3753_/D sky130_fd_sc_hd__a21o_1
Xhold125 _3999_/Q vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _3440_/X vssd1 vssd1 vccd1 vccd1 _3996_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 _3970_/Q vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _3962_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _3382_/X vssd1 vssd1 vccd1 vccd1 _3950_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _3637_/X vssd1 vssd1 vccd1 vccd1 _4079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _3954_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2163__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ _3352_/A _3326_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3326_/X sky130_fd_sc_hd__and3_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3258_/A _3641_/B vssd1 vssd1 vccd1 vccd1 _3257_/Y sky130_fd_sc_hd__nor2_2
X_3188_ _3320_/A _3188_/B vssd1 vssd1 vccd1 vccd1 _3856_/D sky130_fd_sc_hd__or2_1
X_2208_ _2221_/A _2208_/B _2208_/C vssd1 vssd1 vccd1 vccd1 _2208_/X sky130_fd_sc_hd__and3_1
X_2139_ _3933_/Q _3925_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold670 _3856_/Q vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _3850_/Q vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _4084_/Q vssd1 vssd1 vccd1 vccd1 _3646_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2490_ _2332_/X _2487_/Y _2511_/S vssd1 vssd1 vccd1 vccd1 _2491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2145__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3111_ _2988_/B _3102_/D _3157_/A vssd1 vssd1 vccd1 vccd1 _3111_/Y sky130_fd_sc_hd__a21oi_1
X_4091_ _4092_/CLK _4091_/D vssd1 vssd1 vccd1 vccd1 _4091_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3645__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3042_ _3850_/Q _3849_/Q _3851_/Q vssd1 vssd1 vccd1 vccd1 _3043_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ _4089_/CLK _3944_/D vssd1 vssd1 vccd1 vccd1 _3944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2081__B1 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3875_ _4014_/CLK _3875_/D vssd1 vssd1 vccd1 vccd1 _3875_/Q sky130_fd_sc_hd__dfxtp_1
X_2826_ _2667_/X _2815_/X _2825_/X vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3538__A _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2757_ _2674_/X _2742_/X _2756_/X vssd1 vssd1 vccd1 vccd1 _3746_/D sky130_fd_sc_hd__a21o_1
X_2688_ _2688_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _2688_/X sky130_fd_sc_hd__or2_1
XANTENNA__2588__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _2988_/B _3306_/X _3308_/Y vssd1 vssd1 vccd1 vccd1 _3309_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout64 hold700/X vssd1 vssd1 vccd1 vccd1 _3199_/B sky130_fd_sc_hd__clkbuf_8
Xfanout75 _1867_/Y vssd1 vssd1 vccd1 vccd1 _3682_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout86 _3719_/Q vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__buf_4
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout97 _3658_/B vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2127__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1990_ hold580/X _1890_/Y _1989_/X vssd1 vssd1 vccd1 vccd1 _2315_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2063__B1 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3660_ _3506_/A hold269/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3591_ _2619_/A _2613_/Y _3589_/Y _3590_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _3591_/X
+ sky130_fd_sc_hd__o221a_1
X_2611_ _3658_/A _3600_/B vssd1 vssd1 vccd1 vccd1 _3602_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2542_ _3950_/Q hold29/A _3701_/Q _4079_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2543_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2473_ _3947_/Q _3892_/Q _3698_/Q _4076_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2474_/B sky130_fd_sc_hd__mux4_2
X_4074_ _4080_/CLK _4074_/D vssd1 vssd1 vccd1 vccd1 _4074_/Q sky130_fd_sc_hd__dfxtp_1
X_3025_ _3024_/B _3024_/C _3024_/A vssd1 vssd1 vccd1 vccd1 _3056_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3927_ _3938_/CLK _3927_/D vssd1 vssd1 vccd1 vccd1 _3927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3858_ _4029_/CLK _3858_/D vssd1 vssd1 vccd1 vccd1 _3858_/Q sky130_fd_sc_hd__dfxtp_1
X_3789_ _3794_/CLK _3789_/D vssd1 vssd1 vccd1 vccd1 _3789_/Q sky130_fd_sc_hd__dfxtp_1
X_2809_ _2869_/A _2809_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__and3_1
XANTENNA__2357__B2 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2357__A1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2109__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout62_A _2160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1973_ hold93/A _3838_/Q vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3712_ _3795_/CLK _3712_/D vssd1 vssd1 vccd1 vccd1 _3712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3643_ _2655_/X _3640_/X _3642_/X vssd1 vssd1 vccd1 vccd1 _4082_/D sky130_fd_sc_hd__a21o_1
X_3574_ _2630_/A _2646_/D _3573_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _3574_/X sky130_fd_sc_hd__o211a_1
X_2525_ _2524_/X input11/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__mux2_1
X_2456_ _2484_/A _2456_/B vssd1 vssd1 vccd1 vccd1 _2549_/B sky130_fd_sc_hd__or2_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3551__A _3551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2387_ _2677_/A _2551_/B vssd1 vssd1 vccd1 vccd1 _2387_/Y sky130_fd_sc_hd__nand2_1
X_4057_ _4073_/CLK _4057_/D vssd1 vssd1 vccd1 vccd1 _4057_/Q sky130_fd_sc_hd__dfxtp_1
X_3008_ _3065_/B _3008_/B vssd1 vssd1 vccd1 vccd1 _3008_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3463__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3400__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2219_/Y _2287_/X _2308_/Y vssd1 vssd1 vccd1 vccd1 _2310_/Y sky130_fd_sc_hd__a21oi_1
X_3290_ input6/X _1934_/A _3292_/S vssd1 vssd1 vccd1 vccd1 _3290_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2741__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2256_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _2241_/X sky130_fd_sc_hd__or2_1
X_2172_ _2646_/B _2268_/A _2378_/B vssd1 vssd1 vccd1 vccd1 _2172_/X sky130_fd_sc_hd__and3_1
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1956_ _2296_/B _1956_/B vssd1 vssd1 vccd1 vccd1 _1957_/A sky130_fd_sc_hd__or2_1
X_1887_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1887_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout112_A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3626_ _3635_/A0 hold209/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3557_ _3558_/A _3558_/B vssd1 vssd1 vccd1 vccd1 _3559_/A sky130_fd_sc_hd__or2_1
X_2508_ _2508_/A _2508_/B _2508_/C vssd1 vssd1 vccd1 vccd1 _2508_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _3488_/A _3496_/S vssd1 vssd1 vccd1 vccd1 _3488_/Y sky130_fd_sc_hd__nand2_1
X_2439_ _2392_/X _2426_/X _2391_/X vssd1 vssd1 vccd1 vccd1 _2439_/Y sky130_fd_sc_hd__a21oi_1
X_4109_ _4111_/CLK _4109_/D vssd1 vssd1 vccd1 vccd1 _4109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2582__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2790_ _2667_/X _2779_/X _2789_/X vssd1 vssd1 vccd1 vccd1 _3760_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold307 _2933_/X vssd1 vssd1 vccd1 vccd1 _3807_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold329 _3671_/X vssd1 vssd1 vccd1 vccd1 _4102_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _3634_/A0 hold267/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3411_/X sky130_fd_sc_hd__mux2_1
Xhold318 _3877_/Q vssd1 vssd1 vccd1 vccd1 _3222_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2714__B2 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3342_ _3352_/A _3342_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3342_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3656_/A _3273_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3273_/X sky130_fd_sc_hd__and3_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2191_/B _2191_/C _2194_/A vssd1 vssd1 vccd1 vccd1 _2224_/X sky130_fd_sc_hd__a21o_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2151_/X _2154_/X _2155_/S vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__mux2_1
X_2086_ _2222_/A _2208_/B _2208_/C vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__and3_1
XANTENNA__2650__B1 _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2988_ _3157_/A _2988_/B vssd1 vssd1 vccd1 vccd1 _3004_/A sky130_fd_sc_hd__nor2_2
X_1939_ _2616_/A _2616_/C vssd1 vssd1 vccd1 vccd1 _2306_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2180__A _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3609_ _3636_/A0 hold63/X _3612_/S vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2705__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3186__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2944__A1 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _4113_/CLK _3960_/D vssd1 vssd1 vccd1 vccd1 _3960_/Q sky130_fd_sc_hd__dfxtp_1
X_2911_ _3571_/A _3488_/A _1852_/Y hold652/X vssd1 vssd1 vccd1 vccd1 _2911_/X sky130_fd_sc_hd__o22a_1
X_3891_ _4080_/CLK _3891_/D vssd1 vssd1 vccd1 vccd1 _3891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2842_ _2661_/X _2835_/Y _2841_/X vssd1 vssd1 vccd1 vccd1 _3782_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2773_ _2869_/A _2773_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__and3_1
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold126 _3443_/X vssd1 vssd1 vccd1 vccd1 _3999_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _3998_/Q vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _3410_/X vssd1 vssd1 vccd1 vccd1 _3970_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _3400_/X vssd1 vssd1 vccd1 vccd1 _3962_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _3978_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _4050_/Q vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3325_ _2655_/X _3322_/X _3324_/X vssd1 vssd1 vccd1 vccd1 _3325_/X sky130_fd_sc_hd__a21o_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3639_/A0 hold133/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__mux2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2194_/A _2130_/X _2166_/X _2194_/Y _2238_/C vssd1 vssd1 vccd1 vccd1 _2207_/X
+ sky130_fd_sc_hd__a32o_1
X_3187_ hold615/X hold670/X _3189_/S vssd1 vssd1 vccd1 vccd1 _3187_/X sky130_fd_sc_hd__mux2_1
X_2138_ _4086_/Q _3941_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__mux2_1
X_2069_ _3742_/Q _3758_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold660 _3173_/X vssd1 vssd1 vccd1 vccd1 _3174_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _3187_/X vssd1 vssd1 vccd1 vccd1 _3188_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout92_A _3467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3351__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 _4085_/Q vssd1 vssd1 vccd1 vccd1 _3648_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _3175_/X vssd1 vssd1 vccd1 vccd1 _3176_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2813__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2090__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3590__A1 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ _3004_/A _3107_/X _3109_/X _3103_/X _2957_/Y vssd1 vssd1 vccd1 vccd1 _3113_/S
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ _4105_/CLK _4090_/D vssd1 vssd1 vccd1 vccd1 _4090_/Q sky130_fd_sc_hd__dfxtp_1
X_3041_ _3054_/A _3041_/B vssd1 vssd1 vccd1 vccd1 _3051_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ _4088_/CLK _3943_/D vssd1 vssd1 vccd1 vccd1 _3943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2081__A1 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3874_ _4072_/CLK _3874_/D vssd1 vssd1 vccd1 vccd1 _3874_/Q sky130_fd_sc_hd__dfxtp_2
X_2825_ _2863_/A _2825_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2825_/X sky130_fd_sc_hd__and3_1
XFILLER_0_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2756_ _2813_/A _2756_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__and3_1
XANTENNA__3554__A _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2687_ hold688/X _2681_/Y _2686_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3719_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2384__A2 _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3333__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3308_/A _3314_/S vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2519__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3239_ _3247_/A _3239_/B vssd1 vssd1 vccd1 vccd1 _3885_/D sky130_fd_sc_hd__or2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout65 _3554_/A vssd1 vssd1 vccd1 vccd1 _2573_/S sky130_fd_sc_hd__buf_6
Xfanout98 input23/X vssd1 vssd1 vccd1 vccd1 _3658_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout87 _2584_/S1 vssd1 vssd1 vccd1 vccd1 _2582_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout76 _1866_/Y vssd1 vssd1 vccd1 vccd1 _3637_/A0 sky130_fd_sc_hd__buf_4
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3464__A _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 _3779_/Q vssd1 vssd1 vccd1 vccd1 _2831_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3403__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2019__S _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2063__A1 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _3518_/A _3589_/A _2615_/B vssd1 vssd1 vccd1 vccd1 _3590_/X sky130_fd_sc_hd__a21o_1
X_2610_ _2610_/A _2737_/C _2610_/C vssd1 vssd1 vccd1 vccd1 _2733_/S sky130_fd_sc_hd__and3_2
X_2541_ _2564_/A _2541_/B vssd1 vssd1 vccd1 vccd1 _2541_/Y sky130_fd_sc_hd__nand2b_1
X_2472_ _2585_/A _2472_/B vssd1 vssd1 vccd1 vccd1 _2472_/Y sky130_fd_sc_hd__nand2b_1
X_4073_ _4073_/CLK _4073_/D vssd1 vssd1 vccd1 vccd1 _4073_/Q sky130_fd_sc_hd__dfxtp_1
X_3024_ _3024_/A _3024_/B _3024_/C vssd1 vssd1 vccd1 vccd1 _3056_/C sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3690_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3926_ _3938_/CLK _3926_/D vssd1 vssd1 vccd1 vccd1 _3926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3251__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3857_ _3860_/CLK _3857_/D vssd1 vssd1 vccd1 vccd1 _3857_/Q sky130_fd_sc_hd__dfxtp_1
X_2808_ _2667_/X _2797_/X _2807_/X vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__a21o_1
X_3788_ _3794_/CLK _3788_/D vssd1 vssd1 vccd1 vccd1 _3788_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2739_ _2177_/Y _2291_/B _2179_/B vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2045__A1 _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1972_ hold93/A _3838_/Q vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3711_ _3795_/CLK _3711_/D vssd1 vssd1 vccd1 vccd1 _3711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3642_ _3656_/A _3642_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3642_/X sky130_fd_sc_hd__and3_1
XANTENNA__3536__A1 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3573_ _4039_/Q _3579_/B vssd1 vssd1 vccd1 vccd1 _3573_/X sky130_fd_sc_hd__or2_1
X_2524_ _1883_/Y _2523_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__mux2_1
X_2455_ _2372_/Y _2378_/X _2484_/A vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__mux2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ _2318_/X _2337_/Y _2366_/X _2385_/Y vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3551__B _3551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4056_ _4072_/CLK _4056_/D vssd1 vssd1 vccd1 vccd1 _4056_/Q sky130_fd_sc_hd__dfxtp_1
X_3007_ _3106_/A _3004_/Y _3006_/X _3320_/A vssd1 vssd1 vccd1 vccd1 _3007_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2027__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3909_ _4105_/CLK _3909_/D vssd1 vssd1 vccd1 vccd1 _3909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3527__A1 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2122__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2032__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2087_/X _2189_/A _2239_/X vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__a21o_1
X_2171_ _2421_/A _2327_/B vssd1 vssd1 vccd1 vccd1 _2378_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1955_ _3906_/Q _1996_/S _2296_/C _1947_/A vssd1 vssd1 vccd1 vccd1 _1956_/B sky130_fd_sc_hd__o31a_1
XANTENNA__2731__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1886_ _1886_/A vssd1 vssd1 vccd1 vccd1 _1886_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3625_ _1863_/Y hold127/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3625_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout105_A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3556_ _1843_/A _3564_/B _3555_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _4035_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2507_ _2570_/A _2507_/B vssd1 vssd1 vccd1 vccd1 _2508_/C sky130_fd_sc_hd__nand2b_1
X_3487_ _3587_/A _3487_/B vssd1 vssd1 vccd1 vccd1 _4024_/D sky130_fd_sc_hd__and2_1
X_2438_ _2392_/A _2434_/X _2437_/X _2612_/B vssd1 vssd1 vccd1 vccd1 _2438_/X sky130_fd_sc_hd__o211a_1
X_2369_ _2369_/A _2369_/B vssd1 vssd1 vccd1 vccd1 _2484_/A sky130_fd_sc_hd__nand2_2
X_4108_ _4112_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
X_4039_ _4042_/CLK _4039_/D vssd1 vssd1 vccd1 vccd1 _4039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2117__S _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2582__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold308 _3690_/Q vssd1 vssd1 vccd1 vccd1 _3460_/A sky130_fd_sc_hd__buf_2
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3410_ _3633_/A0 hold103/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3410_/X sky130_fd_sc_hd__mux2_1
Xhold319 _3223_/X vssd1 vssd1 vccd1 vccd1 _3877_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3341_ _3341_/A _3641_/A _3640_/C vssd1 vssd1 vccd1 vccd1 _3356_/C sky130_fd_sc_hd__or3b_4
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _2674_/X _3257_/Y _3271_/X vssd1 vssd1 vccd1 vccd1 _3904_/D sky130_fd_sc_hd__a21o_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2222_/B _2187_/X _1995_/Y vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__a21o_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _2152_/X _2153_/X _2160_/A vssd1 vssd1 vccd1 vccd1 _2154_/X sky130_fd_sc_hd__mux2_1
X_2085_ _3693_/Q _2048_/S _2084_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2208_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2650__A1 _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2987_ _2986_/A _2972_/Y _2985_/X _2986_/Y _3131_/A vssd1 vssd1 vccd1 vccd1 _2987_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1938_ _2181_/A _2180_/B vssd1 vssd1 vccd1 vccd1 _1941_/B sky130_fd_sc_hd__nor2_2
XANTENNA__2953__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1869_ _3275_/A vssd1 vssd1 vccd1 vccd1 _3099_/A sky130_fd_sc_hd__inv_2
XANTENNA__2180__B _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3608_ _3635_/A0 hold71/X _3612_/S vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__mux2_1
X_3539_ _3539_/A _3539_/B vssd1 vssd1 vccd1 vccd1 _3539_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3418__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3467__A _3467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2944__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3406__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2880__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3409__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ hold694/X _1853_/Y _1854_/Y _3575_/A _2909_/X vssd1 vssd1 vccd1 vccd1 _2910_/X
+ sky130_fd_sc_hd__o221a_1
X_3890_ _4080_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2841_ _3269_/A _2841_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__and3_1
X_2772_ _2667_/X _2761_/X _2771_/X vssd1 vssd1 vccd1 vccd1 _3752_/D sky130_fd_sc_hd__a21o_1
Xhold105 _3977_/Q vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _3442_/X vssd1 vssd1 vccd1 vccd1 _3998_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _3605_/X vssd1 vssd1 vccd1 vccd1 _4050_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _4063_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _4068_/Q vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2699__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3654_/A _3324_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3324_/X sky130_fd_sc_hd__and3_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3682_/A0 hold119/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__mux2_1
X_2206_ _3654_/B _2306_/B vssd1 vssd1 vccd1 vccd1 _2307_/B sky130_fd_sc_hd__or2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3320_/A _3186_/B vssd1 vssd1 vccd1 vccd1 _3855_/D sky130_fd_sc_hd__or2_1
X_2137_ _2133_/X _2136_/X _2155_/S vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__mux2_1
X_2068_ hold25/A _3798_/Q _2153_/S vssd1 vssd1 vccd1 vccd1 _2068_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold661 _3909_/Q vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _4089_/Q vssd1 vssd1 vccd1 vccd1 _3656_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _3688_/Q vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _4041_/Q vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _3906_/Q vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3639__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2311__B1 _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2862__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2473__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _3040_/A _3040_/B vssd1 vssd1 vccd1 vccd1 _3047_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _4088_/CLK _3942_/D vssd1 vssd1 vccd1 vccd1 _3942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3873_ _4014_/CLK _3873_/D vssd1 vssd1 vccd1 vccd1 _3873_/Q sky130_fd_sc_hd__dfxtp_2
X_2824_ _2664_/X _2815_/X _2823_/X vssd1 vssd1 vccd1 vccd1 _3775_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2755_ _2671_/X _2742_/X _2754_/X vssd1 vssd1 vccd1 vccd1 _3745_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2686_ _2686_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _3136_/A _3307_/B _3307_/C vssd1 vssd1 vccd1 vccd1 _3314_/S sky130_fd_sc_hd__and3b_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2519__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3238_ _1841_/A _3885_/Q _3496_/S vssd1 vssd1 vccd1 vccd1 _3238_/X sky130_fd_sc_hd__mux2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _3275_/C _3169_/B vssd1 vssd1 vccd1 vccd1 _3294_/B sky130_fd_sc_hd__nor2_2
XANTENNA__2844__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout77 _1865_/Y vssd1 vssd1 vccd1 vccd1 _3636_/A0 sky130_fd_sc_hd__buf_4
Xfanout66 _2232_/S vssd1 vssd1 vccd1 vccd1 _3554_/A sky130_fd_sc_hd__clkbuf_8
Xfanout99 _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__buf_4
Xfanout88 _3718_/Q vssd1 vssd1 vccd1 vccd1 _2584_/S1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__2125__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 _3575_/X vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _2832_/X vssd1 vssd1 vccd1 vccd1 _3779_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2599__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3260__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2035__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2446__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2540_ hold85/A _4111_/Q _3966_/Q _3958_/Q _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2541_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2471_ hold91/A hold27/A hold51/A hold11/A _2584_/S0 _3718_/Q vssd1 vssd1 vccd1 vccd1
+ _2472_/B sky130_fd_sc_hd__mux4_1
X_4072_ _4072_/CLK _4072_/D vssd1 vssd1 vccd1 vccd1 _4072_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2826__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3023_ _3191_/A _3027_/A vssd1 vssd1 vccd1 vccd1 _3024_/C sky130_fd_sc_hd__nor2_1
X_3925_ _3938_/CLK _3925_/D vssd1 vssd1 vccd1 vccd1 _3925_/Q sky130_fd_sc_hd__dfxtp_1
X_3856_ _3860_/CLK _3856_/D vssd1 vssd1 vccd1 vccd1 _3856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2807_ _2863_/A _2807_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__and3_1
X_3787_ _3905_/CLK _3787_/D vssd1 vssd1 vccd1 vccd1 _3787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2738_ _2887_/A _2738_/B vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__and2_1
X_2669_ _3656_/A _2669_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2669_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2808__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3710_ _3902_/CLK _3710_/D vssd1 vssd1 vccd1 vccd1 _3710_/Q sky130_fd_sc_hd__dfxtp_1
X_1971_ _3602_/A _1974_/B vssd1 vssd1 vccd1 vccd1 _2940_/A sky130_fd_sc_hd__and2_2
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _3641_/A _3641_/B _3640_/C vssd1 vssd1 vccd1 vccd1 _3656_/C sky130_fd_sc_hd__or3b_2
X_3572_ _2624_/A hold368/X _3571_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _3572_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2523_ _3720_/Q _2520_/Y _2522_/Y _2516_/Y _2518_/Y vssd1 vssd1 vccd1 vccd1 _2523_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2454_ _2571_/B _2454_/B vssd1 vssd1 vccd1 vccd1 _2454_/Y sky130_fd_sc_hd__nor2_1
X_2385_ _2385_/A _2511_/S vssd1 vssd1 vccd1 vccd1 _2385_/Y sky130_fd_sc_hd__nand2_1
Xinput1 custom_settings[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
X_4055_ _4081_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3006_ _2988_/B _2990_/X _3004_/B _3199_/B _2990_/D vssd1 vssd1 vccd1 vccd1 _3006_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3908_ _4105_/CLK _3908_/D vssd1 vssd1 vccd1 vccd1 _3908_/Q sky130_fd_sc_hd__dfxtp_1
X_3839_ _3846_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3215__A1 _3458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _2087_/X _2094_/Y _2169_/X vssd1 vssd1 vccd1 vccd1 _2170_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3206__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1954_ _3321_/B vssd1 vssd1 vccd1 vccd1 _1954_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1885_ _1885_/A vssd1 vssd1 vccd1 vccd1 _1885_/Y sky130_fd_sc_hd__inv_2
X_3624_ _1862_/Y hold187/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3624_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3390__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3555_ _2720_/A _3554_/B _3553_/Y _3554_/Y hold368/X vssd1 vssd1 vccd1 vccd1 _3555_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2193__A1 _3693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2506_ hold638/X _2493_/Y _2505_/X _2492_/X _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3691_/D
+ sky130_fd_sc_hd__o221a_1
X_3486_ _1841_/A hold615/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3487_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2437_ _2435_/X _2436_/X _2512_/A vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__a21o_1
X_2368_ _2646_/B _2119_/S _2319_/X vssd1 vssd1 vccd1 vccd1 _2570_/A sky130_fd_sc_hd__o21ai_4
X_4107_ _4113_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
X_2299_ _2710_/B _2376_/C _2362_/S vssd1 vssd1 vccd1 vccd1 _2571_/A sky130_fd_sc_hd__mux2_4
X_4038_ _4042_/CLK _4038_/D vssd1 vssd1 vccd1 vccd1 _4038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2133__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3381__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2184__A1 _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3684__A1 hold559/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2947__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2043__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 _3221_/X vssd1 vssd1 vccd1 vccd1 _3876_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3340_ _3340_/A _3640_/A _3640_/C vssd1 vssd1 vccd1 vccd1 _3340_/X sky130_fd_sc_hd__and3_2
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__D _3813_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3656_/A _3271_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3271_/X sky130_fd_sc_hd__and3_1
X_2222_ _2222_/A _2222_/B _2222_/C vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__and3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _3778_/Q _3794_/Q _2153_/S vssd1 vssd1 vccd1 vccd1 _2153_/X sky130_fd_sc_hd__mux2_1
X_2084_ _2256_/A _2165_/B _3518_/B vssd1 vssd1 vccd1 vccd1 _2084_/X sky130_fd_sc_hd__and3_1
XFILLER_0_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2986_ _2986_/A _2986_/B vssd1 vssd1 vccd1 vccd1 _2986_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1937_ _3518_/A _2119_/S _2230_/A vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__mux2_4
X_1868_ _3695_/Q vssd1 vssd1 vccd1 vccd1 _1868_/Y sky130_fd_sc_hd__inv_2
X_3607_ _3634_/A0 hold161/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3607_/X sky130_fd_sc_hd__mux2_1
X_3538_ _3540_/A _3538_/B vssd1 vssd1 vccd1 vccd1 _3539_/B sky130_fd_sc_hd__xnor2_1
X_3469_ hold277/X _3470_/B _3468_/Y _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3469_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4112_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3657__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2038__S _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2840_ _2658_/X _2835_/Y _2839_/X vssd1 vssd1 vccd1 vccd1 _3781_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2771_ _2805_/A _2771_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold106 _3418_/X vssd1 vssd1 vccd1 vccd1 _3977_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _4078_/Q vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _4076_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2148__A1 _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold128 _3625_/X vssd1 vssd1 vccd1 vccd1 _4068_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3323_/A _3641_/A _3640_/C vssd1 vssd1 vccd1 vccd1 _3338_/C sky130_fd_sc_hd__or3b_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3637_/A0 hold29/X _3256_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
X_2205_ _3654_/B _2306_/B vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__and2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _4023_/Q hold590/X _3189_/S vssd1 vssd1 vccd1 vccd1 _3185_/X sky130_fd_sc_hd__mux2_1
X_2136_ _2134_/X _2135_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__mux2_1
X_2067_ _3692_/Q _2048_/S _2066_/X _2194_/B vssd1 vssd1 vccd1 vccd1 _2208_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2969_ _3823_/Q _2969_/B vssd1 vssd1 vccd1 vccd1 _3075_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2411__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 _4021_/Q vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 _3914_/Q vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold662 _3283_/X vssd1 vssd1 vccd1 vccd1 _3284_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _4086_/Q vssd1 vssd1 vccd1 vccd1 _3650_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _3494_/X vssd1 vssd1 vccd1 vccd1 _3495_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _3917_/Q vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2473__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3941_ _4088_/CLK _3941_/D vssd1 vssd1 vccd1 vccd1 _3941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3872_ _4072_/CLK _3872_/D vssd1 vssd1 vccd1 vccd1 _3872_/Q sky130_fd_sc_hd__dfxtp_2
X_2823_ _2863_/A _2823_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2823_/X sky130_fd_sc_hd__and3_1
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2754_ _2813_/A _2754_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2754_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2685_ hold520/X _2681_/Y _2684_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ hold640/X _3125_/Y _3303_/X _3305_/X vssd1 vssd1 vccd1 vccd1 _3306_/X sky130_fd_sc_hd__a211o_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3247_/A _3237_/B vssd1 vssd1 vccd1 vccd1 _3884_/D sky130_fd_sc_hd__or2_1
X_3168_ hold302/X _3165_/B _3167_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3168_/X sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2119_ _2115_/X _2118_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2119_/X sky130_fd_sc_hd__mux2_1
X_3099_ _3099_/A _3833_/Q _3099_/C vssd1 vssd1 vccd1 vccd1 _3100_/C sky130_fd_sc_hd__or3_1
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout78 _1864_/Y vssd1 vssd1 vccd1 vccd1 _3635_/A0 sky130_fd_sc_hd__buf_4
Xfanout89 _2584_/S0 vssd1 vssd1 vccd1 vccd1 _2582_/S0 sky130_fd_sc_hd__buf_6
Xfanout67 _2159_/S vssd1 vssd1 vccd1 vccd1 _2152_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2930__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2141__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold470 _3754_/Q vssd1 vssd1 vccd1 vccd1 _2775_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _3755_/Q vssd1 vssd1 vccd1 vccd1 _2777_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _3710_/Q vssd1 vssd1 vccd1 vccd1 _2657_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2446__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2470_ _2585_/A _2469_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2470_/Y sky130_fd_sc_hd__a21oi_1
X_4071_ _4072_/CLK _4071_/D vssd1 vssd1 vccd1 vccd1 _4071_/Q sky130_fd_sc_hd__dfxtp_1
X_3022_ hold597/X _3020_/Y _3021_/X vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3924_ _3938_/CLK _3924_/D vssd1 vssd1 vccd1 vccd1 _3924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3855_ _3860_/CLK _3855_/D vssd1 vssd1 vccd1 vccd1 _3855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2806_ _2664_/X _2797_/X _2805_/X vssd1 vssd1 vccd1 vccd1 _3767_/D sky130_fd_sc_hd__a21o_1
X_3786_ _3902_/CLK _3786_/D vssd1 vssd1 vccd1 vccd1 _3786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3795_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2737_ _2737_/A _2737_/B _2737_/C vssd1 vssd1 vccd1 vccd1 _2740_/S sky130_fd_sc_hd__and3_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2668_ _2652_/Y _2667_/X _2666_/X vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2599_ _3635_/A0 hold255/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2599_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2136__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2753__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1970_ _2230_/A _2158_/S _1959_/C _1959_/D _1969_/X vssd1 vssd1 vccd1 vccd1 _1974_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ _3640_/A _3640_/B _3640_/C vssd1 vssd1 vccd1 vccd1 _3640_/X sky130_fd_sc_hd__and3_2
XFILLER_0_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3571_ _3571_/A _3579_/B vssd1 vssd1 vccd1 vccd1 _3571_/X sky130_fd_sc_hd__or2_1
X_2522_ _2585_/A _2522_/B vssd1 vssd1 vccd1 vccd1 _2522_/Y sky130_fd_sc_hd__nand2_1
X_2453_ _2334_/Y _2335_/X _2304_/Y vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__a21oi_1
X_2384_ _2573_/S _2296_/B _1942_/B _2256_/A vssd1 vssd1 vccd1 vccd1 _2551_/B sky130_fd_sc_hd__a31o_2
X_4123_ _4123_/A vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__buf_1
Xinput2 custom_settings[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4054_ _4073_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
X_3005_ _3118_/B _3001_/X _3004_/Y _3114_/A vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_78_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3907_ _4105_/CLK _3907_/D vssd1 vssd1 vccd1 vccd1 _3907_/Q sky130_fd_sc_hd__dfxtp_1
X_3838_ _3862_/CLK _3838_/D vssd1 vssd1 vccd1 vccd1 _3838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3769_ _3794_/CLK _3769_/D vssd1 vssd1 vccd1 vccd1 _3769_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout60_A _2155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1953_ _1959_/D _3529_/A _2646_/B vssd1 vssd1 vccd1 vccd1 _3321_/B sky130_fd_sc_hd__mux2_4
XANTENNA__2504__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1884_ _1884_/A vssd1 vssd1 vccd1 vccd1 _1884_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3623_ _3676_/A0 hold219/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3623_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2717__B2 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ _3554_/A _3554_/B vssd1 vssd1 vccd1 vccd1 _3554_/Y sky130_fd_sc_hd__nor2_1
X_2505_ _2393_/B _2504_/X _2493_/Y vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__a21bo_1
X_3485_ _3497_/A _3485_/B vssd1 vssd1 vccd1 vccd1 _4023_/D sky130_fd_sc_hd__and2_1
X_2436_ _2418_/X _2432_/Y _2551_/B vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__a21o_1
X_2367_ _2318_/X _2337_/Y _2366_/X vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__a21o_1
X_4106_ _4111_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
X_2298_ _2710_/B _2296_/X _2297_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2376_/C sky130_fd_sc_hd__o22a_1
X_4037_ _4042_/CLK _4037_/D vssd1 vssd1 vccd1 vccd1 _4037_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2956__A1 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2500__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2947__A1 hold536/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1922__A2 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3270_ _2671_/X _3257_/Y _3269_/X vssd1 vssd1 vccd1 vccd1 _3903_/D sky130_fd_sc_hd__a21o_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2221_/A _2221_/B _2221_/C vssd1 vssd1 vccd1 vccd1 _2221_/X sky130_fd_sc_hd__and3_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _3770_/Q _3754_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2152_/X sky130_fd_sc_hd__mux2_1
X_2083_ _2074_/X _2082_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3518_/B sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2985_ _2974_/B _2984_/Y _3818_/Q vssd1 vssd1 vccd1 vccd1 _2985_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ _4100_/Q _1890_/Y _1934_/X vssd1 vssd1 vccd1 vccd1 _2155_/S sky130_fd_sc_hd__o21a_4
X_1867_ _3694_/Q vssd1 vssd1 vccd1 vccd1 _1867_/Y sky130_fd_sc_hd__inv_2
X_3606_ _3633_/A0 hold151/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3606_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3573__B _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3537_ _3529_/A _3529_/B _3536_/X vssd1 vssd1 vccd1 vccd1 _3538_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3363__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3468_ _3468_/A _3470_/B vssd1 vssd1 vccd1 vccd1 _3468_/Y sky130_fd_sc_hd__nand2_1
X_3399_ _3676_/A0 hold185/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3399_/X sky130_fd_sc_hd__mux2_1
X_2419_ _2229_/B _2373_/B _2424_/B vssd1 vssd1 vccd1 vccd1 _2420_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3290__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3658__B _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2054__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2770_ _2664_/X _2761_/X _2769_/X vssd1 vssd1 vccd1 vccd1 _3751_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold107 _3986_/Q vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _4113_/Q vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3345__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold118 _3636_/X vssd1 vssd1 vccd1 vccd1 _4078_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1906__B _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3322_/A _3640_/A _3640_/C vssd1 vssd1 vccd1 vccd1 _3322_/X sky130_fd_sc_hd__and3_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3636_/A0 hold17/X _3256_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
X_3184_ _3320_/A _3184_/B vssd1 vssd1 vccd1 vccd1 _3854_/D sky130_fd_sc_hd__or2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _3544_/S _2203_/X _2606_/B vssd1 vssd1 vccd1 vccd1 _2306_/B sky130_fd_sc_hd__a21oi_1
X_2135_ _3776_/Q _3792_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2135_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2066_ _2256_/A _2165_/B _3525_/B vssd1 vssd1 vccd1 vccd1 _2066_/X sky130_fd_sc_hd__and3_1
XANTENNA__3281__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2968_ _3150_/B _2968_/B vssd1 vssd1 vccd1 vccd1 _3157_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1919_ _1919_/A _1919_/B vssd1 vssd1 vccd1 vccd1 _1919_/Y sky130_fd_sc_hd__nand2_1
X_2899_ _3140_/B _2899_/B _3140_/C vssd1 vssd1 vccd1 vccd1 _3088_/A sky130_fd_sc_hd__or3_1
Xhold630 _3879_/Q vssd1 vssd1 vccd1 vccd1 _1860_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold652 _4042_/Q vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _3852_/Q vssd1 vssd1 vccd1 vccd1 _3179_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold663 _4049_/Q vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 _3818_/Q vssd1 vssd1 vccd1 vccd1 _2976_/B sky130_fd_sc_hd__buf_1
Xhold685 _3824_/Q vssd1 vssd1 vccd1 vccd1 _2997_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _3301_/X vssd1 vssd1 vccd1 vccd1 _3302_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2928__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3327__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3940_ _4088_/CLK _3940_/D vssd1 vssd1 vccd1 vccd1 _3940_/Q sky130_fd_sc_hd__dfxtp_1
X_3871_ _4072_/CLK _3871_/D vssd1 vssd1 vccd1 vccd1 _3871_/Q sky130_fd_sc_hd__dfxtp_1
X_2822_ _2661_/X _2815_/X _2821_/X vssd1 vssd1 vccd1 vccd1 _3774_/D sky130_fd_sc_hd__a21o_1
X_2753_ _2667_/X _2742_/X _2752_/X vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2684_ _2684_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _4025_/Q _3124_/Y _3304_/Y _4017_/Q vssd1 vssd1 vccd1 vccd1 _3305_/X sky130_fd_sc_hd__a22o_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3564_/A _3884_/Q _3494_/S vssd1 vssd1 vccd1 vccd1 _3236_/X sky130_fd_sc_hd__mux2_1
X_3167_ _3846_/Q _3157_/A _3148_/A _3154_/Y vssd1 vssd1 vccd1 vccd1 _3167_/X sky130_fd_sc_hd__a211o_1
X_3098_ _3123_/B _3125_/A _3095_/X _3097_/A vssd1 vssd1 vccd1 vccd1 _3115_/B sky130_fd_sc_hd__o211a_1
X_2118_ _2116_/X _2117_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3254__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2049_ _2192_/A _2220_/B _2031_/X vssd1 vssd1 vccd1 vccd1 _2049_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout79 _1863_/Y vssd1 vssd1 vccd1 vccd1 _3634_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout57 _3494_/S vssd1 vssd1 vccd1 vccd1 _3496_/S sky130_fd_sc_hd__clkbuf_8
Xfanout68 _2153_/S vssd1 vssd1 vccd1 vccd1 _2159_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 _3941_/Q vssd1 vssd1 vccd1 vccd1 _3368_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 _3774_/Q vssd1 vssd1 vccd1 vccd1 _2821_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _2778_/X vssd1 vssd1 vccd1 vccd1 _3755_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _3904_/Q vssd1 vssd1 vccd1 vccd1 _3271_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2048__A1 _3695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3548__A1 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4073_/CLK _4070_/D vssd1 vssd1 vccd1 vccd1 _4070_/Q sky130_fd_sc_hd__dfxtp_1
X_3021_ _3861_/Q _3050_/C _3020_/Y hold597/X vssd1 vssd1 vccd1 vccd1 _3021_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3923_ _3939_/CLK _3923_/D vssd1 vssd1 vccd1 vccd1 _3923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3854_ _3860_/CLK _3854_/D vssd1 vssd1 vccd1 vccd1 _3854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2805_ _2805_/A _2805_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3785_ _3902_/CLK _3785_/D vssd1 vssd1 vccd1 vccd1 _3785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2736_ _2887_/A _2736_/B vssd1 vssd1 vccd1 vccd1 _3738_/D sky130_fd_sc_hd__and2_1
X_2667_ _2332_/X _2489_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2598_ _3634_/A0 hold189/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2278__A1 _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ _3691_/Q _2681_/Y _3218_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3219_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2202__A1 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold290 _4012_/Q vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _1841_/A _3564_/B _3569_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _4037_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2062__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2521_ _3949_/Q hold17/A _3700_/Q _4078_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2522_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2452_ _3458_/A _2439_/Y _2451_/X _2438_/X _2698_/A vssd1 vssd1 vccd1 vccd1 _3689_/D
+ sky130_fd_sc_hd__o221a_1
X_2383_ _2573_/S _2296_/B _1942_/B _2256_/A vssd1 vssd1 vccd1 vccd1 _2511_/S sky130_fd_sc_hd__a31oi_4
X_4122_ _4123_/A vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__buf_1
X_4053_ _4081_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
Xinput3 io_in[10] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_3004_ _3004_/A _3004_/B vssd1 vssd1 vccd1 vccd1 _3004_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2761__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3906_ _4105_/CLK _3906_/D vssd1 vssd1 vccd1 vccd1 _3906_/Q sky130_fd_sc_hd__dfxtp_1
X_3837_ _4077_/CLK _3837_/D vssd1 vssd1 vccd1 vccd1 _3837_/Q sky130_fd_sc_hd__dfxtp_1
X_3768_ _3791_/CLK _3768_/D vssd1 vssd1 vccd1 vccd1 _3768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ hold35/X _2708_/Y _2741_/S _2678_/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__a22o_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3699_ _4080_/CLK _3699_/D vssd1 vssd1 vccd1 vccd1 _3699_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3448__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3620__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3439__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1952_ hold673/X hold312/X _1996_/S vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__mux2_8
XANTENNA__3611__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1883_ _1883_/A vssd1 vssd1 vccd1 vccd1 _1883_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3622_ _3874_/Q _3873_/Q _3675_/B vssd1 vssd1 vccd1 vccd1 _3630_/S sky130_fd_sc_hd__or3_4
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3553_ _3553_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3553_/Y sky130_fd_sc_hd__xnor2_1
X_2504_ _2503_/X input12/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__mux2_1
X_3484_ _3564_/A hold669/X _3494_/S vssd1 vssd1 vccd1 vccd1 _3485_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3678__A0 _1863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2435_ _2435_/A _2511_/S vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2366_ _2508_/A _2508_/B vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__and2_1
X_4105_ _4105_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__2756__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2297_ _3554_/A _1942_/B _2737_/C _2610_/A vssd1 vssd1 vccd1 vccd1 _2297_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ _4101_/CLK _4036_/D vssd1 vssd1 vccd1 vccd1 _4036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2500__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2956__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3669__A0 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2947__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2220_/A _2220_/B vssd1 vssd1 vccd1 vccd1 _2220_/X sky130_fd_sc_hd__or2_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2151_ _2149_/X _2150_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2151_/X sky130_fd_sc_hd__mux2_1
X_2082_ _1959_/C _2077_/X _2079_/X _2081_/X vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2635__A1 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2984_ _3820_/Q _2984_/B vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__nand2_1
X_1935_ hold592/X _1890_/Y _1934_/X vssd1 vssd1 vccd1 vccd1 _1959_/C sky130_fd_sc_hd__o21ai_4
XANTENNA__2494__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1866_ _3693_/Q vssd1 vssd1 vccd1 vccd1 _1866_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3605_ _3676_/A0 hold137/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout103_A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ _3529_/A _3529_/B _3531_/B vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__o21ba_1
X_3467_ _3467_/A _3467_/B vssd1 vssd1 vccd1 vccd1 _4014_/D sky130_fd_sc_hd__or2_1
X_2418_ _2571_/B _2415_/X _2417_/Y _2508_/A vssd1 vssd1 vccd1 vccd1 _2418_/X sky130_fd_sc_hd__a211o_1
X_3398_ _3675_/A _3613_/C vssd1 vssd1 vccd1 vccd1 _3406_/S sky130_fd_sc_hd__or2_4
X_2349_ _3518_/A _2349_/B vssd1 vssd1 vccd1 vccd1 _2349_/X sky130_fd_sc_hd__and2_1
XANTENNA__2874__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4019_ _4092_/CLK _4019_/D vssd1 vssd1 vccd1 vccd1 _4019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2396__A _2592_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold108 _3429_/X vssd1 vssd1 vccd1 vccd1 _3986_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2070__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold119 _3896_/Q vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_3321_ _3321_/A _3321_/B vssd1 vssd1 vccd1 vccd1 _3640_/C sky130_fd_sc_hd__nor2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3635_/A0 hold13/X _3256_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
X_3183_ hold645/X hold677/X _3189_/S vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2856__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2227_/S _3558_/A _2197_/Y _2279_/S vssd1 vssd1 vccd1 vccd1 _2203_/X sky130_fd_sc_hd__o2bb2a_1
X_2134_ _3768_/Q _3752_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2134_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2737__C _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2065_ _2056_/X _2064_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3525_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3939_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2967_ _2967_/A _3824_/Q _3163_/A _2997_/C vssd1 vssd1 vccd1 vccd1 _2968_/B sky130_fd_sc_hd__and4_1
XANTENNA__2467__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2898_ _3134_/B _3163_/A _3134_/C vssd1 vssd1 vccd1 vccd1 _2988_/B sky130_fd_sc_hd__and3_4
X_1918_ _1919_/A _1919_/B vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__and2_1
X_1849_ _4025_/Q vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__inv_2
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold620 _3501_/X vssd1 vssd1 vccd1 vccd1 _4030_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _3859_/Q vssd1 vssd1 vccd1 vccd1 _3193_/A sky130_fd_sc_hd__buf_1
Xhold631 _3226_/X vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 _3180_/X vssd1 vssd1 vccd1 vccd1 _3852_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _2590_/X vssd1 vssd1 vccd1 vccd1 _3695_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _2975_/X vssd1 vssd1 vccd1 vccd1 _2977_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _2997_/Y vssd1 vssd1 vccd1 vccd1 _2998_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _3830_/Q vssd1 vssd1 vccd1 vccd1 _3100_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3519_ _3507_/A _2277_/B _3502_/X _3502_/B _3506_/A vssd1 vssd1 vccd1 vccd1 _3520_/B
+ sky130_fd_sc_hd__a32oi_2
XANTENNA__3272__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2155__S _2155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2480__C1 _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2838__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _4105_/CLK _3870_/D vssd1 vssd1 vccd1 vccd1 _3870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2821_ _2863_/A _2821_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2821_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2752_ _2805_/A _2752_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2752_/X sky130_fd_sc_hd__and3_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2683_ hold559/X _2681_/Y _2682_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__o211a_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _3304_/A _3304_/B vssd1 vssd1 vccd1 vccd1 _3304_/Y sky130_fd_sc_hd__nor2_1
X_3235_ _3497_/A _3235_/B vssd1 vssd1 vccd1 vccd1 _3883_/D sky130_fd_sc_hd__nand2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3148_/A _3164_/X hold380/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__o211a_1
X_3097_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3097_/Y sky130_fd_sc_hd__inv_2
X_2117_ _3777_/Q _3793_/Q _2153_/S vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3579__B _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2048_ _2277_/B _3695_/Q _2048_/S vssd1 vssd1 vccd1 vccd1 _2220_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3999_ _4014_/CLK _3999_/D vssd1 vssd1 vccd1 vccd1 _3999_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout58 _2937_/X vssd1 vssd1 vccd1 vccd1 _3494_/S sky130_fd_sc_hd__buf_4
Xfanout69 _2153_/S vssd1 vssd1 vccd1 vccd1 _2161_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold461 _3926_/Q vssd1 vssd1 vccd1 vccd1 _3334_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _3751_/Q vssd1 vssd1 vccd1 vccd1 _2769_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _3795_/Q vssd1 vssd1 vccd1 vccd1 _2869_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _3792_/Q vssd1 vssd1 vccd1 vccd1 _2863_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _3728_/Q vssd1 vssd1 vccd1 vccd1 _2706_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020_ _3193_/A _3024_/B vssd1 vssd1 vccd1 vccd1 _3020_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3922_ _3939_/CLK _3922_/D vssd1 vssd1 vccd1 vccd1 _3922_/Q sky130_fd_sc_hd__dfxtp_1
X_3853_ _4029_/CLK _3853_/D vssd1 vssd1 vccd1 vccd1 _3853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2804_ _2661_/X _2797_/X _2803_/X vssd1 vssd1 vccd1 vccd1 _3766_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3784_ _3902_/CLK _3784_/D vssd1 vssd1 vccd1 vccd1 _3784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2735_ _2732_/A _2734_/X _2735_/S vssd1 vssd1 vccd1 vccd1 _2736_/B sky130_fd_sc_hd__mux2_1
X_2666_ _3269_/A _2666_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__and3_1
XANTENNA__3172__B1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2597_ _3633_/A0 hold217/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4031_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3218_ _3218_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _3218_/X sky130_fd_sc_hd__or2_1
X_3149_ hold288/X _3165_/B _3148_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold280 _3458_/Y vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _3463_/X vssd1 vssd1 vccd1 vccd1 _4012_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3466__A1 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2520_ _2585_/A _2520_/B vssd1 vssd1 vccd1 vccd1 _2520_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2451_ _2393_/B _2450_/X _2439_/Y vssd1 vssd1 vccd1 vccd1 _2451_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2382_ _2367_/X _2385_/A _2381_/Y vssd1 vssd1 vccd1 vccd1 _2382_/Y sky130_fd_sc_hd__a21oi_1
X_4052_ _4073_/CLK _4052_/D vssd1 vssd1 vccd1 vccd1 _4052_/Q sky130_fd_sc_hd__dfxtp_1
Xinput4 io_in[16] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _3118_/B _3120_/A _3163_/B vssd1 vssd1 vccd1 vccd1 _3004_/B sky130_fd_sc_hd__and3_1
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3209__A1 _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3905_ _3905_/CLK _3905_/D vssd1 vssd1 vccd1 vccd1 _3905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3836_ _4095_/CLK _3836_/D vssd1 vssd1 vccd1 vccd1 _3836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3767_ _3767_/CLK _3767_/D vssd1 vssd1 vccd1 vccd1 _3767_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3393__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2718_ hold7/X _2708_/Y _2741_/S _2674_/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__a22o_1
X_3698_ _4095_/CLK _3698_/D vssd1 vssd1 vccd1 vccd1 _3698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2649_ _2296_/B _2737_/B _2677_/B vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2671__A2 _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3384__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2662__A2 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1951_ hold563/X _1890_/Y _1949_/X vssd1 vssd1 vccd1 vccd1 _2164_/S sky130_fd_sc_hd__o21ai_4
X_1882_ _1882_/A vssd1 vssd1 vccd1 vccd1 _1882_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2073__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3621_ _3639_/A0 hold145/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ _3550_/Y _3552_/B vssd1 vssd1 vccd1 vccd1 _3553_/B sky130_fd_sc_hd__and2b_1
X_2503_ _1884_/Y _2502_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__mux2_1
X_3483_ _3587_/A _3483_/B vssd1 vssd1 vccd1 vccd1 _4022_/D sky130_fd_sc_hd__and2_1
X_2434_ _2573_/S _2433_/X _3558_/B vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__a21o_1
X_2365_ _2348_/Y _2454_/B _2571_/B vssd1 vssd1 vccd1 vccd1 _2508_/B sky130_fd_sc_hd__mux2_1
X_4104_ _4105_/CLK _4104_/D vssd1 vssd1 vccd1 vccd1 _4104_/Q sky130_fd_sc_hd__dfxtp_1
X_2296_ _3544_/S _2296_/B _2296_/C vssd1 vssd1 vccd1 vccd1 _2296_/X sky130_fd_sc_hd__or3_1
X_4035_ _4042_/CLK _4035_/D vssd1 vssd1 vccd1 vccd1 _4035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3819_ _3860_/CLK _3819_/D vssd1 vssd1 vccd1 vccd1 _3819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2158__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _3746_/Q _3762_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2068__S _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2081_ _2158_/S _2080_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__o21a_1
X_2983_ _3131_/A _2983_/B _2983_/C vssd1 vssd1 vccd1 vccd1 _2983_/X sky130_fd_sc_hd__and3_1
XFILLER_0_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1934_ _1934_/A _1996_/S vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__or2_2
XFILLER_0_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2494__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1865_ _3692_/Q vssd1 vssd1 vccd1 vccd1 _1865_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3604_ _3874_/Q _3873_/Q _3604_/C vssd1 vssd1 vccd1 vccd1 _3612_/S sky130_fd_sc_hd__or3_4
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3535_ _1845_/A _3564_/B _3533_/Y _3534_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _4033_/D
+ sky130_fd_sc_hd__o221a_1
X_3466_ hold347/X _3637_/A0 _3470_/B vssd1 vssd1 vccd1 vccd1 _3466_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2417_ _2571_/A _2333_/Y _2416_/Y _2571_/B vssd1 vssd1 vccd1 vccd1 _2417_/Y sky130_fd_sc_hd__a211oi_1
X_3397_ _3871_/Q _3454_/A _3872_/Q vssd1 vssd1 vccd1 vccd1 _3613_/C sky130_fd_sc_hd__or3b_2
X_2348_ _2550_/B vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__inv_2
X_2279_ _3507_/B _3498_/B _2279_/S vssd1 vssd1 vccd1 vccd1 _2280_/B sky130_fd_sc_hd__mux2_1
X_4018_ _4031_/CLK _4018_/D vssd1 vssd1 vccd1 vccd1 _4018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold109 _4005_/Q vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2553__A1 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3320_ _3320_/A _3320_/B vssd1 vssd1 vccd1 vccd1 _3920_/D sky130_fd_sc_hd__or2_1
XFILLER_0_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3634_/A0 hold177/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__mux2_1
X_3182_ _3247_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _3853_/D sky130_fd_sc_hd__or2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _3633_/A0 _2646_/B _2197_/Y _2201_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2606_/B
+ sky130_fd_sc_hd__o221a_1
X_2133_ _2131_/X _2132_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2133_/X sky130_fd_sc_hd__mux2_1
X_2064_ _1959_/C _2059_/X _2061_/X _2063_/X vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2966_ _2964_/X _2965_/X _3163_/A vssd1 vssd1 vccd1 vccd1 _3150_/B sky130_fd_sc_hd__o21a_1
XANTENNA__2467__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2897_ _2960_/A _3824_/Q vssd1 vssd1 vccd1 vccd1 _3140_/C sky130_fd_sc_hd__or2_1
X_1917_ _3602_/A _3600_/B hold286/X vssd1 vssd1 vccd1 vccd1 _1919_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1848_ _4030_/Q vssd1 vssd1 vccd1 vccd1 _1848_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2792__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold621 _4047_/Q vssd1 vssd1 vccd1 vccd1 _2621_/A sky130_fd_sc_hd__buf_1
Xhold610 _3687_/X vssd1 vssd1 vccd1 vccd1 _3874_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold654 _3194_/X vssd1 vssd1 vccd1 vccd1 _3859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 _3816_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 hold742/X vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold687 _2998_/X vssd1 vssd1 vccd1 vccd1 _3824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _4031_/Q vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold676 _3100_/Y vssd1 vssd1 vccd1 vccd1 _3294_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _3518_/A _3518_/B vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__xnor2_1
X_3449_ _3635_/A0 hold43/X _3453_/S vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__mux2_1
Xhold698 _2977_/X vssd1 vssd1 vccd1 vccd1 _3818_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ _2658_/X _2815_/X _2819_/X vssd1 vssd1 vccd1 vccd1 _2820_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2751_ _2664_/X _2742_/X _2750_/X vssd1 vssd1 vccd1 vccd1 _3743_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2774__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2682_ _2682_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _2682_/X sky130_fd_sc_hd__or2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _3050_/A _3832_/Q _2923_/B _3084_/Y vssd1 vssd1 vccd1 vccd1 _3303_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3234_ _1843_/Y _1856_/Y _3496_/S vssd1 vssd1 vccd1 vccd1 _3234_/X sky130_fd_sc_hd__mux2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3165_/A _3165_/B vssd1 vssd1 vccd1 vccd1 _3165_/X sky130_fd_sc_hd__or2_1
X_3096_ _3830_/Q _3829_/Q _3099_/C _3132_/B vssd1 vssd1 vccd1 vccd1 _3097_/A sky130_fd_sc_hd__or4_1
X_2116_ _3769_/Q _3753_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__mux2_1
X_2047_ _2045_/Y _2046_/Y _2164_/S _2038_/X vssd1 vssd1 vccd1 vccd1 _2277_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2462__B1 _3551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3998_ _4014_/CLK _3998_/D vssd1 vssd1 vccd1 vccd1 _3998_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2780__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout59 _1988_/Y vssd1 vssd1 vccd1 vccd1 _3554_/B sky130_fd_sc_hd__buf_4
X_2949_ hold547/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold451 _3940_/Q vssd1 vssd1 vccd1 vccd1 _3366_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 _3898_/Q vssd1 vssd1 vccd1 vccd1 _3259_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2939__B _2939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 _3782_/Q vssd1 vssd1 vccd1 vccd1 _2841_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _2864_/X vssd1 vssd1 vccd1 vccd1 _3792_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _3769_/Q vssd1 vssd1 vccd1 vccd1 _2809_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _2870_/X vssd1 vssd1 vccd1 vccd1 _3795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4095_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3469__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3921_ _3939_/CLK _3921_/D vssd1 vssd1 vccd1 vccd1 _3921_/Q sky130_fd_sc_hd__dfxtp_1
X_3852_ _4029_/CLK _3852_/D vssd1 vssd1 vccd1 vccd1 _3852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2803_ _2805_/A _2803_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__and3_1
XANTENNA__2747__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3783_ _3902_/CLK _3783_/D vssd1 vssd1 vccd1 vccd1 _3783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2734_ _2378_/A _2733_/X _2734_/S vssd1 vssd1 vccd1 vccd1 _2734_/X sky130_fd_sc_hd__mux2_1
X_2665_ _2652_/Y _2664_/X _2663_/X vssd1 vssd1 vccd1 vccd1 _3712_/D sky130_fd_sc_hd__a21o_1
X_2596_ _3676_/A0 hold253/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1970__A2 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3217_ _3688_/Q _3201_/Y _3216_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3217_/X sky130_fd_sc_hd__o211a_1
X_3148_ _3148_/A _3148_/B vssd1 vssd1 vccd1 vccd1 _3148_/X sky130_fd_sc_hd__or2_1
X_3079_ _3120_/C _2989_/B _3078_/X _3077_/X _2899_/B vssd1 vssd1 vccd1 vccd1 _3080_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 _3660_/X vssd1 vssd1 vccd1 vccd1 _4091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _3459_/X vssd1 vssd1 vccd1 vccd1 _4010_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _3843_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2521__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2450_ _2449_/X input14/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2381_ hold672/X _2385_/A _2573_/S vssd1 vssd1 vccd1 vccd1 _2381_/Y sky130_fd_sc_hd__o21ai_1
X_4051_ _4073_/CLK _4051_/D vssd1 vssd1 vccd1 vccd1 _4051_/Q sky130_fd_sc_hd__dfxtp_1
Xinput5 io_in[17] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_3002_ _3004_/A _2990_/X hold578/X _3001_/X _3320_/A vssd1 vssd1 vccd1 vccd1 _3002_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1939__A _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3904_ _3905_/CLK _3904_/D vssd1 vssd1 vccd1 vccd1 _3904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3835_ _4077_/CLK _3835_/D vssd1 vssd1 vccd1 vccd1 _3835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3766_ _3791_/CLK _3766_/D vssd1 vssd1 vccd1 vccd1 _3766_/Q sky130_fd_sc_hd__dfxtp_1
X_2717_ hold87/X _2708_/Y _2741_/S _2671_/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__a22o_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3697_ _4080_/CLK _3697_/D vssd1 vssd1 vccd1 vccd1 _3697_/Q sky130_fd_sc_hd__dfxtp_1
X_2648_ _2677_/B vssd1 vssd1 vccd1 vccd1 _2648_/Y sky130_fd_sc_hd__inv_2
X_2579_ _2585_/A _2579_/B vssd1 vssd1 vccd1 vccd1 _2579_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ hold563/X _1890_/Y _1949_/X vssd1 vssd1 vccd1 vccd1 _1959_/D sky130_fd_sc_hd__o21a_2
X_1881_ _1881_/A vssd1 vssd1 vccd1 vccd1 _1881_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _3682_/A0 hold233/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3620_/X sky130_fd_sc_hd__mux2_1
X_3551_ _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3552_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3375__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2502_ _3720_/Q _2499_/Y _2501_/Y _2495_/Y _2497_/Y vssd1 vssd1 vccd1 vccd1 _2502_/X
+ sky130_fd_sc_hd__a32o_1
X_3482_ _1843_/A hold645/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2433_ _3458_/A _2426_/X _2432_/Y _2418_/X vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__a22o_1
X_2364_ _2347_/S _2416_/B _2363_/X vssd1 vssd1 vccd1 vccd1 _2454_/B sky130_fd_sc_hd__o21ai_1
X_4103_ _4103_/CLK _4103_/D vssd1 vssd1 vccd1 vccd1 _4103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2295_ _1941_/B _2178_/B _2293_/Y _2349_/B vssd1 vssd1 vccd1 vccd1 _2295_/X sky130_fd_sc_hd__a211o_1
X_4034_ _4042_/CLK _4034_/D vssd1 vssd1 vccd1 vccd1 _4034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3818_ _3860_/CLK _3818_/D vssd1 vssd1 vccd1 vccd1 _3818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3749_ _3791_/CLK _3749_/D vssd1 vssd1 vccd1 vccd1 _3749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3357__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ _3900_/Q _3782_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2080_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2873__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2982_ _2982_/A _2982_/B vssd1 vssd1 vccd1 vccd1 _2986_/B sky130_fd_sc_hd__nand2_1
X_1933_ hold611/X hold257/X _1996_/S vssd1 vssd1 vccd1 vccd1 _3518_/A sky130_fd_sc_hd__mux2_8
X_1864_ _3691_/Q vssd1 vssd1 vccd1 vccd1 _1864_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3603_ _2614_/B _3602_/Y _3467_/A vssd1 vssd1 vccd1 vccd1 _4049_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3534_ _3592_/A _3554_/B hold368/X vssd1 vssd1 vccd1 vccd1 _3534_/X sky130_fd_sc_hd__a21o_1
X_3465_ hold275/X _3470_/B _3464_/Y _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3465_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2416_ _2571_/A _2416_/B vssd1 vssd1 vccd1 vccd1 _2416_/Y sky130_fd_sc_hd__nor2_1
X_3396_ _3639_/A0 hold131/X _3396_/S vssd1 vssd1 vccd1 vccd1 _3396_/X sky130_fd_sc_hd__mux2_1
X_2347_ _2427_/B _2571_/D _2347_/S vssd1 vssd1 vccd1 vccd1 _2550_/B sky130_fd_sc_hd__mux2_1
X_2278_ _3544_/S _3507_/B _2277_/X vssd1 vssd1 vccd1 vccd1 _3498_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _4031_/CLK _4017_/D vssd1 vssd1 vccd1 vccd1 _4017_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2007__B _2232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3339__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1862__A _3458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2677__B _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3633_/A0 hold247/X _3256_/S vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__mux2_1
X_3181_ _4021_/Q hold553/X _3189_/S vssd1 vssd1 vccd1 vccd1 _3181_/X sky130_fd_sc_hd__mux2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2378_/A _2424_/A _2424_/B _2230_/A vssd1 vssd1 vccd1 vccd1 _2201_/X sky130_fd_sc_hd__a211o_1
X_2132_ _3744_/Q _3760_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2132_/X sky130_fd_sc_hd__mux2_1
X_2063_ _2158_/S _2062_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2063_/X sky130_fd_sc_hd__o21a_1
X_2965_ _3140_/B _3120_/C _2997_/C _3076_/B vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__a2bb2o_1
X_2896_ _2960_/A _3824_/Q vssd1 vssd1 vccd1 vccd1 _3134_/C sky130_fd_sc_hd__nor2_1
X_1916_ _2008_/C _3600_/B _3910_/Q vssd1 vssd1 vccd1 vccd1 _1919_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1847_ _4031_/Q vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3767_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 _3007_/Y vssd1 vssd1 vccd1 vccd1 _3828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _3916_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold633 _3236_/X vssd1 vssd1 vccd1 vccd1 _3237_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _2956_/Y vssd1 vssd1 vccd1 vccd1 _3816_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 _3599_/X vssd1 vssd1 vccd1 vccd1 _4047_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3517_ _3517_/A _3517_/B vssd1 vssd1 vccd1 vccd1 _3517_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold677 _3854_/Q vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _3512_/X vssd1 vssd1 vccd1 vccd1 _4031_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 _3913_/Q vssd1 vssd1 vccd1 vccd1 _1949_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _3693_/Q vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__buf_1
X_3448_ _3634_/A0 hold9/X _3453_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
Xhold699 _3817_/Q vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
X_3379_ _3634_/A0 hold163/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3379_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2480__A1 _3460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3420__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2750_ _2805_/A _2750_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2681_ _3201_/A _2681_/B vssd1 vssd1 vccd1 vccd1 _2681_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _3601_/A _3302_/B vssd1 vssd1 vccd1 vccd1 _3917_/D sky130_fd_sc_hd__and2_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3497_/A _3233_/B vssd1 vssd1 vccd1 vccd1 _3882_/D sky130_fd_sc_hd__nand2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ hold294/X _3199_/B _3157_/X _3163_/X vssd1 vssd1 vccd1 vccd1 _3164_/X sky130_fd_sc_hd__o22a_1
X_3095_ _3834_/Q _3833_/Q _3829_/Q _3832_/Q vssd1 vssd1 vccd1 vccd1 _3095_/X sky130_fd_sc_hd__or4b_1
X_2115_ _2113_/X _2114_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2046_ _1959_/C _2041_/X _1959_/D vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__a21oi_1
X_3997_ _4016_/CLK _3997_/D vssd1 vssd1 vccd1 vccd1 _3997_/Q sky130_fd_sc_hd__dfxtp_1
X_2948_ _3636_/A0 _2940_/X _2947_/Y vssd1 vssd1 vccd1 vccd1 _2948_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3411__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2879_ _2887_/A _2879_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__and3_1
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold463 _3799_/Q vssd1 vssd1 vccd1 vccd1 _2879_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _3740_/Q vssd1 vssd1 vccd1 vccd1 _2744_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _3796_/Q vssd1 vssd1 vccd1 vccd1 _2873_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _3260_/X vssd1 vssd1 vccd1 vccd1 _3898_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _3933_/Q vssd1 vssd1 vccd1 vccd1 _3350_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _3768_/Q vssd1 vssd1 vccd1 vccd1 _2807_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _3902_/Q vssd1 vssd1 vccd1 vccd1 _3267_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold368_A _2646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout69_A _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3402__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2881__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _4095_/CLK _3920_/D vssd1 vssd1 vccd1 vccd1 _3920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3851_ _4029_/CLK _3851_/D vssd1 vssd1 vccd1 vccd1 _3851_/Q sky130_fd_sc_hd__dfxtp_1
X_2802_ _2658_/X _2797_/X _2801_/X vssd1 vssd1 vccd1 vccd1 _2802_/X sky130_fd_sc_hd__a21o_1
X_3782_ _3902_/CLK _3782_/D vssd1 vssd1 vccd1 vccd1 _3782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2733_ _2732_/X _3566_/A _2733_/S vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2664_ _2361_/X _2510_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__mux2_8
X_2595_ _3871_/Q _3631_/A _3872_/Q vssd1 vssd1 vccd1 vccd1 _2603_/S sky130_fd_sc_hd__or3b_4
XANTENNA__1970__A3 _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3216_ _1889_/Y _3201_/A _2410_/B _2408_/A vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__a31o_1
X_3147_ hold271/X _2989_/B _3199_/B vssd1 vssd1 vccd1 vccd1 _3148_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2683__A1 hold559/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3078_ _3106_/A _3118_/B _3120_/A vssd1 vssd1 vccd1 vccd1 _3078_/X sky130_fd_sc_hd__or3_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2791__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3632__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2029_ _2256_/A _2165_/B _3682_/A0 vssd1 vssd1 vccd1 vccd1 _2192_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold271 _3840_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _3618_/X vssd1 vssd1 vccd1 vccd1 _4062_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _4016_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _3156_/X vssd1 vssd1 vccd1 vccd1 _3843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3623__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2521__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1937__A0 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3139__C1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2362__A0 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2380_ _2375_/X _2507_/B _2570_/A vssd1 vssd1 vccd1 vccd1 _2385_/A sky130_fd_sc_hd__mux2_2
X_4050_ _4073_/CLK _4050_/D vssd1 vssd1 vccd1 vccd1 _4050_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 io_in[18] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _3120_/A _3163_/B _3004_/A vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__and3_1
XANTENNA__3614__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3903_ _3939_/CLK _3903_/D vssd1 vssd1 vccd1 vccd1 _3903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3834_ _4095_/CLK _3834_/D vssd1 vssd1 vccd1 vccd1 _3834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3765_ _3791_/CLK _3765_/D vssd1 vssd1 vccd1 vccd1 _3765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2716_ hold19/X _2708_/Y _2741_/S _2667_/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__a22o_1
X_3696_ _4080_/CLK _3696_/D vssd1 vssd1 vccd1 vccd1 _3696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2647_ _2647_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2677_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2578_ _3976_/Q _4073_/Q _4065_/Q _4057_/Q _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2579_/B sky130_fd_sc_hd__mux4_1
XANTENNA__2353__B1 _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3605__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1865__A _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2344__B1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2696__A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3320__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ input3/X vssd1 vssd1 vccd1 vccd1 _1880_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3550_/Y sky130_fd_sc_hd__nor2_1
X_2501_ _2564_/A _2501_/B vssd1 vssd1 vccd1 vccd1 _2501_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3481_ _3497_/A _3481_/B vssd1 vssd1 vccd1 vccd1 _4021_/D sky130_fd_sc_hd__and2_1
X_2432_ _2508_/A _2431_/Y _2426_/X vssd1 vssd1 vccd1 vccd1 _2432_/Y sky130_fd_sc_hd__a21oi_1
X_2363_ _2362_/S _2355_/Y _2349_/X _2571_/A vssd1 vssd1 vccd1 vccd1 _2363_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2886__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4102_ _4105_/CLK _4102_/D vssd1 vssd1 vccd1 vccd1 _4102_/Q sky130_fd_sc_hd__dfxtp_1
X_4033_ _4042_/CLK _4033_/D vssd1 vssd1 vccd1 vccd1 _4033_/Q sky130_fd_sc_hd__dfxtp_1
X_2294_ _1941_/B _2178_/B _2293_/Y vssd1 vssd1 vccd1 vccd1 _2677_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3599__C1 _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2810__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3817_ _3862_/CLK _3817_/D vssd1 vssd1 vccd1 vccd1 _3817_/Q sky130_fd_sc_hd__dfxtp_2
X_3748_ _3795_/CLK _3748_/D vssd1 vssd1 vccd1 vccd1 _3748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ _1864_/Y hold213/X _3683_/S vssd1 vssd1 vccd1 vccd1 _3679_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2868__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3315__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output32_A _2939_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2592__C _2592_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2981_ _2982_/A _2982_/B vssd1 vssd1 vccd1 vccd1 _2983_/B sky130_fd_sc_hd__or2_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1932_ _2230_/A _3554_/A _2227_/S vssd1 vssd1 vccd1 vccd1 _2296_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1863_ _3460_/A vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__inv_2
Xinput20 io_in[7] vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__clkbuf_1
X_3602_ _3602_/A _3602_/B vssd1 vssd1 vccd1 vccd1 _3602_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3533_ _3554_/B _3533_/B vssd1 vssd1 vccd1 vccd1 _3533_/Y sky130_fd_sc_hd__nor2_1
X_3464_ _3692_/Q _3470_/B vssd1 vssd1 vccd1 vccd1 _3464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2415_ _2571_/A _2314_/X _2316_/X _2414_/Y vssd1 vssd1 vccd1 vccd1 _2415_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3395_ _3682_/A0 hold15/X _3396_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
XANTENNA__2403__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2346_ _3507_/A _2345_/X _2362_/S vssd1 vssd1 vccd1 vccd1 _2571_/D sky130_fd_sc_hd__mux2_1
X_2277_ _3554_/A _2277_/B vssd1 vssd1 vccd1 vccd1 _2277_/X sky130_fd_sc_hd__or2_1
X_4016_ _4016_/CLK _4016_/D vssd1 vssd1 vccd1 vccd1 _4016_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2492__C1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3578__A2 _2646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2230_/A _2424_/B vssd1 vssd1 vccd1 vccd1 _2200_/Y sky130_fd_sc_hd__nor2_1
X_3180_ hold637/X _3189_/S _3179_/X _3497_/A vssd1 vssd1 vccd1 vccd1 _3180_/X sky130_fd_sc_hd__o211a_1
X_2131_ hold19/A _3800_/Q _2153_/S vssd1 vssd1 vccd1 vccd1 _2131_/X sky130_fd_sc_hd__mux2_1
X_2062_ _3901_/Q _3783_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2062_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2095__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3266__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2964_ _3823_/Q _2969_/B _3076_/B _2961_/X vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__a31o_1
X_1915_ _3507_/A vssd1 vssd1 vccd1 vccd1 _3581_/A sky130_fd_sc_hd__inv_2
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2895_ _2990_/D _3118_/B _3120_/A vssd1 vssd1 vccd1 vccd1 _2899_/B sky130_fd_sc_hd__or3_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1846_ _1846_/A vssd1 vssd1 vccd1 vccd1 _1846_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2124__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 _3299_/X vssd1 vssd1 vccd1 vccd1 _3300_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold601 _3827_/Q vssd1 vssd1 vccd1 vccd1 _3118_/B sky130_fd_sc_hd__buf_2
Xhold645 _4022_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__buf_1
Xhold623 _3835_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
X_3516_ _3506_/A _3506_/B _3506_/X _3507_/X vssd1 vssd1 vccd1 vccd1 _3517_/B sky130_fd_sc_hd__a22oi_2
XANTENNA_fanout101_A _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 _3907_/Q vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 _4088_/Q vssd1 vssd1 vccd1 vccd1 _3654_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _3183_/X vssd1 vssd1 vccd1 vccd1 _3184_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 _3292_/X vssd1 vssd1 vccd1 vccd1 _3293_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3447_ _3633_/A0 hold33/X _3453_/S vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__mux2_1
Xhold689 _3686_/X vssd1 vssd1 vccd1 vccd1 _3873_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3378_ _3633_/A0 hold221/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3378_/X sky130_fd_sc_hd__mux2_1
X_2329_ _2246_/Y _2284_/X _2235_/Y vssd1 vssd1 vccd1 vccd1 _2329_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2680_ _3201_/A _2681_/B vssd1 vssd1 vccd1 vccd1 _3224_/B sky130_fd_sc_hd__and2_2
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2879__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3301_ input7/X hold673/X _3301_/S vssd1 vssd1 vccd1 vccd1 _3301_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _1844_/Y _1857_/Y _3494_/S vssd1 vssd1 vccd1 vccd1 _3232_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3163_/A _3163_/B vssd1 vssd1 vccd1 vccd1 _3163_/X sky130_fd_sc_hd__and2_1
X_2114_ _3745_/Q _3761_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ _3829_/Q _3036_/X _3132_/B _3093_/X vssd1 vssd1 vccd1 vccd1 _3102_/B sky130_fd_sc_hd__o211a_1
X_2045_ _2151_/S _2043_/X _2044_/X vssd1 vssd1 vccd1 vccd1 _2045_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3996_ _4016_/CLK _3996_/D vssd1 vssd1 vccd1 vccd1 _3996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ hold536/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2947_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2878_ _2661_/X _2871_/X _2877_/X vssd1 vssd1 vccd1 vccd1 _3798_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold420 _3937_/Q vssd1 vssd1 vccd1 vccd1 _3360_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 _3745_/Q vssd1 vssd1 vccd1 vccd1 _2754_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _2874_/X vssd1 vssd1 vccd1 vccd1 _3796_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _2745_/X vssd1 vssd1 vccd1 vccd1 _3740_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _2808_/X vssd1 vssd1 vccd1 vccd1 _3768_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _3746_/Q vssd1 vssd1 vccd1 vccd1 _2756_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _3786_/Q vssd1 vssd1 vccd1 vccd1 _2849_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 _3777_/Q vssd1 vssd1 vccd1 vccd1 _2827_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__C1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1868__A _3695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _4029_/CLK _3850_/D vssd1 vssd1 vccd1 vccd1 _3850_/Q sky130_fd_sc_hd__dfxtp_1
X_2801_ _2805_/A _2801_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2801_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3781_ _3902_/CLK _3781_/D vssd1 vssd1 vccd1 vccd1 _3781_/Q sky130_fd_sc_hd__dfxtp_1
X_2732_ _2732_/A _2732_/B vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2663_ _2869_/A _2663_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2663_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2594_ _3454_/A _2594_/B vssd1 vssd1 vccd1 vccd1 _3631_/A sky130_fd_sc_hd__or2_2
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3215_ _3458_/A _3201_/Y _3214_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3215_/X sky130_fd_sc_hd__o211a_1
X_3146_ hold271/X _3165_/B _3145_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__o211a_1
X_3077_ _2990_/C _3077_/B _3119_/B vssd1 vssd1 vccd1 vccd1 _3077_/X sky130_fd_sc_hd__and3b_1
X_2028_ _2019_/X _2027_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3502_/B sky130_fd_sc_hd__mux2_2
X_3979_ _4112_/CLK hold92/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3396__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold261 _4073_/Q vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 _3489_/X vssd1 vssd1 vccd1 vccd1 _4025_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold283 _3471_/X vssd1 vssd1 vccd1 vccd1 _4016_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _3146_/X vssd1 vssd1 vccd1 vccd1 _3840_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _3845_/Q vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold478_A _3808_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1937__A1 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_in[19] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3000_ _3163_/B _3004_/A _3120_/A vssd1 vssd1 vccd1 vccd1 _3000_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2665__A2 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3902_ _3902_/CLK _3902_/D vssd1 vssd1 vccd1 vccd1 _3902_/Q sky130_fd_sc_hd__dfxtp_1
X_3833_ _4095_/CLK _3833_/D vssd1 vssd1 vccd1 vccd1 _3833_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3378__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3764_ _3795_/CLK _3764_/D vssd1 vssd1 vccd1 vccd1 _3764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3695_ _4011_/CLK _3695_/D vssd1 vssd1 vccd1 vccd1 _3695_/Q sky130_fd_sc_hd__dfxtp_2
X_2715_ hold31/X _2708_/Y _2741_/S _2664_/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__a22o_1
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2646_ _3467_/A _2646_/B _3554_/A _2646_/D vssd1 vssd1 vccd1 vccd1 _2647_/B sky130_fd_sc_hd__or4_4
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2577_ _2393_/X _2572_/S _2390_/Y vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2656__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3129_ hold302/X hold700/X _3128_/X vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3480_ _1844_/A hold640/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3481_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2500_ _3948_/Q hold13/A _3699_/Q hold57/A _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2501_/B sky130_fd_sc_hd__mux4_2
X_2431_ _2571_/B _2427_/X _2428_/X _2430_/Y vssd1 vssd1 vccd1 vccd1 _2431_/Y sky130_fd_sc_hd__a31oi_2
XANTENNA__2887__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2362_ _3529_/A _2361_/X _2362_/S vssd1 vssd1 vccd1 vccd1 _2416_/B sky130_fd_sc_hd__mux2_1
X_2293_ _2291_/X _2292_/Y _2182_/X vssd1 vssd1 vccd1 vccd1 _2293_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2098__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4101_ _4101_/CLK _4101_/D vssd1 vssd1 vccd1 vccd1 _4101_/Q sky130_fd_sc_hd__dfxtp_1
X_4032_ _4045_/CLK _4032_/D vssd1 vssd1 vccd1 vccd1 _4032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4089_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3816_ _4077_/CLK _3816_/D vssd1 vssd1 vccd1 vccd1 _3816_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3747_ _3778_/CLK _3747_/D vssd1 vssd1 vccd1 vccd1 _3747_/Q sky130_fd_sc_hd__dfxtp_1
X_3678_ _1863_/Y hold27/X _3683_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
X_2629_ _2630_/A _2629_/B vssd1 vssd1 vccd1 vccd1 _2637_/C sky130_fd_sc_hd__and2_1
XFILLER_0_80_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _2984_/B _2978_/B _2979_/Y vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1931_ hold683/X hold328/X _1996_/S vssd1 vssd1 vccd1 vccd1 _2232_/S sky130_fd_sc_hd__mux2_4
X_1862_ _3458_/A vssd1 vssd1 vccd1 vccd1 _1862_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 io_in[24] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
Xinput21 io_in[8] vssd1 vssd1 vccd1 vccd1 _1882_/A sky130_fd_sc_hd__clkbuf_1
X_3601_ _3601_/A _3602_/B _3601_/C vssd1 vssd1 vccd1 vccd1 _4048_/D sky130_fd_sc_hd__and3_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3532_ _3528_/Y _3531_/Y _3554_/A vssd1 vssd1 vccd1 vccd1 _3533_/B sky130_fd_sc_hd__mux2_1
X_3463_ hold290/X _3470_/B _3462_/Y _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3463_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2414_ _2362_/S _2670_/A _2328_/Y _2571_/A vssd1 vssd1 vccd1 vccd1 _2414_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__3506__A _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2410__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3394_ _3637_/A0 hold111/X _3396_/S vssd1 vssd1 vccd1 vccd1 _3394_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2403__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2345_ _2344_/X _2616_/A _2345_/S vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__mux2_1
X_2276_ _2238_/B _2223_/X _2224_/X _2274_/X _2275_/X vssd1 vssd1 vccd1 vccd1 _3507_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4015_ _4016_/CLK _4015_/D vssd1 vssd1 vccd1 vccd1 _4015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2011__A3 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2786__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2397__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2130_ _3690_/Q _2048_/S _2129_/X _2194_/B vssd1 vssd1 vccd1 vccd1 _2130_/X sky130_fd_sc_hd__a211o_1
X_2061_ _2142_/A _2061_/B vssd1 vssd1 vccd1 vccd1 _2061_/X sky130_fd_sc_hd__or2_1
X_2963_ _2967_/A _3824_/Q vssd1 vssd1 vccd1 vccd1 _3076_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ hold651/X hold316/X _1996_/S vssd1 vssd1 vccd1 vccd1 _3507_/A sky130_fd_sc_hd__mux2_8
XFILLER_0_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2894_ _2990_/D _3118_/B _3120_/A vssd1 vssd1 vccd1 vccd1 _3163_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1845_ _1845_/A vssd1 vssd1 vccd1 vccd1 _1845_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold602 _3005_/X vssd1 vssd1 vccd1 vccd1 _3827_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold624 _3091_/X vssd1 vssd1 vccd1 vccd1 _3835_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3513_/Y _3515_/B vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__nand2b_1
Xhold635 _3279_/X vssd1 vssd1 vccd1 vccd1 _3280_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 _3874_/Q vssd1 vssd1 vccd1 vccd1 _2688_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _4026_/Q vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__buf_1
Xhold657 _3918_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 _3737_/Q vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _4082_/Q vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3446_ _1861_/Y hold195/X _3453_/S vssd1 vssd1 vccd1 vccd1 _3446_/X sky130_fd_sc_hd__mux2_1
X_3377_ _3676_/A0 hold239/X _3384_/S vssd1 vssd1 vccd1 vccd1 _3377_/X sky130_fd_sc_hd__mux2_1
X_2328_ _2362_/S _3551_/B vssd1 vssd1 vccd1 vccd1 _2328_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2701__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3846_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2259_ _2604_/B _2261_/C _4084_/Q vssd1 vssd1 vccd1 vccd1 _2350_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2768__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2315__A _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2759__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3300_ _3601_/A _3300_/B vssd1 vssd1 vccd1 vccd1 _3916_/D sky130_fd_sc_hd__and2_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3497_/A _3231_/B vssd1 vssd1 vccd1 vccd1 _3881_/D sky130_fd_sc_hd__nand2_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ hold294/X _3165_/B _3161_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3162_/X sky130_fd_sc_hd__o211a_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ hold87/A _3801_/Q _2153_/S vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__mux2_1
X_3093_ _3832_/Q _3123_/B _3304_/A vssd1 vssd1 vccd1 vccd1 _3093_/X sky130_fd_sc_hd__or3_1
X_2044_ _2142_/A _2042_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2542__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3995_ _4011_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
X_2946_ _3637_/A0 _2940_/X _2945_/Y vssd1 vssd1 vccd1 vccd1 _2946_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2877_ _2887_/A _2877_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__and3_1
Xhold410 _3776_/Q vssd1 vssd1 vccd1 vccd1 _2825_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _3361_/X vssd1 vssd1 vccd1 vccd1 _3937_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold454 _3757_/Q vssd1 vssd1 vccd1 vccd1 _2783_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _3772_/Q vssd1 vssd1 vccd1 vccd1 _2817_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _3903_/Q vssd1 vssd1 vccd1 vccd1 _3269_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _3762_/Q vssd1 vssd1 vccd1 vccd1 _2793_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _3794_/Q vssd1 vssd1 vccd1 vccd1 _2867_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 _3712_/Q vssd1 vssd1 vccd1 vccd1 _2663_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3429_ _3633_/A0 hold107/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3429_/X sky130_fd_sc_hd__mux2_1
Xhold498 _3722_/Q vssd1 vssd1 vccd1 vccd1 _2694_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2800_ _2655_/X _2797_/X _2799_/X vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__a21o_1
X_3780_ _3902_/CLK _3780_/D vssd1 vssd1 vccd1 vccd1 _3780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2601__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2731_ _2887_/A _2731_/B vssd1 vssd1 vccd1 vccd1 _3737_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2662_ _2652_/Y _2661_/X _2660_/X vssd1 vssd1 vccd1 vccd1 _3711_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2593_ _3874_/Q _3873_/Q vssd1 vssd1 vccd1 vccd1 _2594_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3514__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _1889_/Y _3201_/A _2410_/B _2408_/B vssd1 vssd1 vccd1 vccd1 _3214_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3145_ _3199_/B _3144_/X _3148_/A vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__a21o_1
X_3076_ _3134_/B _3076_/B vssd1 vssd1 vccd1 vccd1 _3119_/B sky130_fd_sc_hd__nand2_1
X_2027_ _1959_/C _2022_/X _2024_/X _2026_/X vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2515__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3978_ _4112_/CLK _3978_/D vssd1 vssd1 vccd1 vccd1 _3978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2929_ hold300/X _2925_/Y _2928_/X _3601_/A vssd1 vssd1 vccd1 vccd1 _2929_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1946__A2 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold251 _4110_/Q vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _3630_/X vssd1 vssd1 vccd1 vccd1 _4073_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 _3377_/X vssd1 vssd1 vccd1 vccd1 _3945_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _4011_/Q vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _3162_/X vssd1 vssd1 vccd1 vccd1 _3845_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _3806_/Q vssd1 vssd1 vccd1 vccd1 _1989_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold638_A _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 io_in[22] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output55_A _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_2_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3901_ _3902_/CLK _3901_/D vssd1 vssd1 vccd1 vccd1 _3901_/Q sky130_fd_sc_hd__dfxtp_1
X_3832_ _4092_/CLK _3832_/D vssd1 vssd1 vccd1 vccd1 _3832_/Q sky130_fd_sc_hd__dfxtp_1
X_3763_ _3778_/CLK _3763_/D vssd1 vssd1 vccd1 vccd1 _3763_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1928__A2 _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3694_ _4011_/CLK _3694_/D vssd1 vssd1 vccd1 vccd1 _3694_/Q sky130_fd_sc_hd__dfxtp_1
X_2714_ hold25/X _2708_/Y _2741_/S _2661_/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__a22o_1
X_2645_ _2645_/A _2645_/B vssd1 vssd1 vccd1 vccd1 _3708_/D sky130_fd_sc_hd__nor2_1
X_2576_ _2392_/A _2573_/X _2575_/X _2612_/B vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2271__A1_N _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128_ _2988_/B _3127_/X _3120_/Y _3157_/A vssd1 vssd1 vccd1 vccd1 _3128_/X sky130_fd_sc_hd__a211o_1
X_3059_ _3010_/Y _3058_/X _3114_/A vssd1 vssd1 vccd1 vccd1 _3059_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3369__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3541__A1 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2430_ _2571_/B _2430_/B vssd1 vssd1 vccd1 vccd1 _2430_/Y sky130_fd_sc_hd__nor2_1
X_2361_ _1941_/B _2356_/B _2357_/X _2360_/Y vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__o2bb2a_1
X_4100_ _4101_/CLK _4100_/D vssd1 vssd1 vccd1 vccd1 _4100_/Q sky130_fd_sc_hd__dfxtp_1
X_2292_ _2291_/A _2291_/B _2180_/B vssd1 vssd1 vccd1 vccd1 _2292_/Y sky130_fd_sc_hd__a21oi_1
X_4031_ _4031_/CLK _4031_/D vssd1 vssd1 vccd1 vccd1 _4031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3815_ _4113_/CLK _3815_/D vssd1 vssd1 vccd1 vccd1 _3815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3746_ _3794_/CLK _3746_/D vssd1 vssd1 vccd1 vccd1 _3746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3677_ _1862_/Y hold59/X _3683_/S vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__mux2_1
XANTENNA__1982__A _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2628_ _2624_/A _2640_/B _2627_/Y _3227_/A vssd1 vssd1 vccd1 vccd1 _3704_/D sky130_fd_sc_hd__o211a_1
X_2559_ hold5/A _3999_/Q _4015_/Q hold67/A _2582_/S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1
+ _2559_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3450__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1930_ hold328/X _1996_/S _1929_/Y vssd1 vssd1 vccd1 vccd1 _1930_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2253__B2 _3693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1861_ _3688_/Q vssd1 vssd1 vccd1 vccd1 _1861_/Y sky130_fd_sc_hd__inv_2
Xinput11 io_in[25] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
Xinput22 io_in[9] vssd1 vssd1 vccd1 vccd1 _1881_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3600_ _3658_/A _3600_/B vssd1 vssd1 vccd1 vccd1 _3601_/C sky130_fd_sc_hd__or2_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3531_ _3531_/A _3531_/B vssd1 vssd1 vccd1 vccd1 _3531_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3462_ _3691_/Q _3470_/B vssd1 vssd1 vccd1 vccd1 _3462_/Y sky130_fd_sc_hd__nand2_1
X_3393_ _3636_/A0 hold101/X _3396_/S vssd1 vssd1 vccd1 vccd1 _3393_/X sky130_fd_sc_hd__mux2_1
X_2413_ hold672/X _2394_/X _2412_/X _2389_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3688_/D
+ sky130_fd_sc_hd__o221a_1
X_2344_ _3642_/B _2181_/A _1945_/Y _2280_/B vssd1 vssd1 vccd1 vccd1 _2344_/X sky130_fd_sc_hd__a22o_1
X_2275_ _2220_/A _2220_/B _2093_/B vssd1 vssd1 vccd1 vccd1 _2275_/X sky130_fd_sc_hd__o21a_1
X_4014_ _4014_/CLK _4014_/D vssd1 vssd1 vccd1 vccd1 _4014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3441__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2244__A1 _2232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _4045_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3432__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4081_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2397__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2060_ _3712_/Q _3724_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2061_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3671__A0 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3423__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2962_ _2962_/A _2969_/B vssd1 vssd1 vccd1 vccd1 _2989_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _2369_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _2834_/A sky130_fd_sc_hd__and2_2
X_2893_ _2962_/A _2992_/A vssd1 vssd1 vccd1 vccd1 _3140_/B sky130_fd_sc_hd__or2_2
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1844_ _1844_/A vssd1 vssd1 vccd1 vccd1 _1844_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold603 _3888_/Q vssd1 vssd1 vccd1 vccd1 _1853_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold625 _3915_/Q vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _4094_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _3518_/A _3514_/B vssd1 vssd1 vccd1 vccd1 _3515_/B sky130_fd_sc_hd__nand2_1
Xhold614 _2689_/X vssd1 vssd1 vccd1 vccd1 _3720_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 _4023_/Q vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _3822_/Q vssd1 vssd1 vccd1 vccd1 _2992_/A sky130_fd_sc_hd__clkbuf_2
Xhold658 _3310_/X vssd1 vssd1 vccd1 vccd1 _3918_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3445_ _3445_/A _3455_/A vssd1 vssd1 vccd1 vccd1 _3453_/S sky130_fd_sc_hd__or2_4
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3872_/Q _3871_/Q _3631_/A vssd1 vssd1 vccd1 vccd1 _3384_/S sky130_fd_sc_hd__or3_4
XANTENNA__2162__B1 _2155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2567__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2327_ _3544_/S _2327_/B vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__and2_2
X_2258_ _2604_/B _2261_/C vssd1 vssd1 vccd1 vccd1 _2258_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3662__A0 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2189_ _2189_/A _2189_/B _2189_/C vssd1 vssd1 vccd1 vccd1 _2197_/A sky130_fd_sc_hd__and3_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3414__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2217__A1 _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2477__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3405__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _1845_/Y _1858_/Y _3496_/S vssd1 vssd1 vccd1 vccd1 _3230_/X sky130_fd_sc_hd__mux2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2144__B1 _2155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3161_ _3844_/Q _3157_/A _3148_/A _3154_/Y vssd1 vssd1 vccd1 vccd1 _3161_/X sky130_fd_sc_hd__a211o_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2695__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2112_ _3688_/Q _2048_/S _2111_/X vssd1 vssd1 vccd1 vccd1 _2238_/C sky130_fd_sc_hd__a21o_1
X_3092_ _3099_/A _3833_/Q vssd1 vssd1 vccd1 vccd1 _3132_/B sky130_fd_sc_hd__nand2_1
X_2043_ _3898_/Q _3780_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2043_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2542__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3994_ _4011_/CLK _3994_/D vssd1 vssd1 vccd1 vccd1 _3994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2945_ hold583/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2945_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2876_ _2658_/X _2871_/X _2875_/X vssd1 vssd1 vccd1 vccd1 _3797_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold400 _3758_/Q vssd1 vssd1 vccd1 vccd1 _2785_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _2826_/X vssd1 vssd1 vccd1 vccd1 _3776_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _3942_/Q vssd1 vssd1 vccd1 vccd1 _3370_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold740/X vssd1 vssd1 vccd1 vccd1 _1845_/A sky130_fd_sc_hd__buf_1
Xhold433 _2818_/X vssd1 vssd1 vccd1 vccd1 _3772_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold466 _3924_/Q vssd1 vssd1 vccd1 vccd1 _3330_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _2784_/X vssd1 vssd1 vccd1 vccd1 _3757_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _3725_/Q vssd1 vssd1 vccd1 vccd1 _2700_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3681__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold499 _3810_/Q vssd1 vssd1 vccd1 vccd1 hold499/X sky130_fd_sc_hd__dlygate4sd3_1
X_3428_ _1861_/Y hold49/X _3435_/S vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
Xhold488 _3781_/Q vssd1 vssd1 vccd1 vccd1 _2839_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3641_/A _3359_/B _3640_/C vssd1 vssd1 vccd1 vccd1 _3374_/C sky130_fd_sc_hd__or3b_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3635__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2061__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2126__B1 _2155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2730_ hold679/X _2729_/X _2735_/S vssd1 vssd1 vccd1 vccd1 _2731_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2661_ _2355_/Y _2531_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2592_ _2939_/A _2592_/B _2592_/C _2940_/A vssd1 vssd1 vccd1 vccd1 _3454_/A sky130_fd_sc_hd__or4b_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3213_ _3460_/A _3201_/Y _3212_/X _3687_/C1 vssd1 vssd1 vccd1 vccd1 _3213_/X sky130_fd_sc_hd__o211a_1
X_3144_ _3163_/A _2964_/X _3157_/B vssd1 vssd1 vccd1 vccd1 _3144_/X sky130_fd_sc_hd__a21o_1
X_3075_ _3824_/Q _3075_/B vssd1 vssd1 vccd1 vccd1 _3077_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3617__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2026_ _2158_/S _2025_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2026_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2515__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2840__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3676__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3977_ _4111_/CLK _3977_/D vssd1 vssd1 vccd1 vccd1 _3977_/Q sky130_fd_sc_hd__dfxtp_1
X_2928_ input5/X _3834_/Q _3072_/B vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__or3_1
XFILLER_0_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2863_/A _2859_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__and3_1
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3002__D1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 _3403_/X vssd1 vssd1 vccd1 vccd1 _3965_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _3680_/X vssd1 vssd1 vccd1 vccd1 _4110_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold241 _3700_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _3461_/X vssd1 vssd1 vccd1 vccd1 _4011_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _4058_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _3842_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _2931_/X vssd1 vssd1 vccd1 vccd1 _3806_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2108__B1 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout67_A _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2442__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 io_in[23] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2822__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3900_ _3902_/CLK _3900_/D vssd1 vssd1 vccd1 vccd1 _3900_/Q sky130_fd_sc_hd__dfxtp_1
X_3831_ _4092_/CLK _3831_/D vssd1 vssd1 vccd1 vccd1 _3831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3762_ _3794_/CLK _3762_/D vssd1 vssd1 vccd1 vccd1 _3762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2713_ hold47/X _2708_/Y _2741_/S _2658_/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__a22o_1
X_3693_ _4014_/CLK _3693_/D vssd1 vssd1 vccd1 vccd1 _3693_/Q sky130_fd_sc_hd__dfxtp_2
X_2644_ _2642_/A _2640_/B _3227_/A vssd1 vssd1 vccd1 vccd1 _2645_/B sky130_fd_sc_hd__o21ai_1
X_2575_ _2511_/S _2572_/S _2571_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3525__A _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3127_ _4028_/Q _3088_/B _3095_/X _3126_/X vssd1 vssd1 vccd1 vccd1 _3127_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3058_ _3065_/B _3058_/B vssd1 vssd1 vccd1 vccd1 _3058_/X sky130_fd_sc_hd__and2b_1
X_2009_ _2009_/A _2009_/B _2008_/C vssd1 vssd1 vccd1 vccd1 _2646_/D sky130_fd_sc_hd__or3b_4
XFILLER_0_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2804__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2360_ _2360_/A _2360_/B vssd1 vssd1 vccd1 vccd1 _2360_/Y sky130_fd_sc_hd__nor2_1
X_2291_ _2291_/A _2291_/B vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__or2_1
X_4030_ _4031_/CLK _4030_/D vssd1 vssd1 vccd1 vccd1 _4030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3814_ _4113_/CLK _3814_/D vssd1 vssd1 vccd1 vccd1 _3814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3745_ _3778_/CLK _3745_/D vssd1 vssd1 vccd1 vccd1 _3745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3676_ _3676_/A0 hold55/X _3683_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
XFILLER_0_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2627_ _2640_/B _2627_/B vssd1 vssd1 vccd1 vccd1 _2627_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4047_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2558_ _2564_/A _2558_/B vssd1 vssd1 vccd1 vccd1 _2558_/Y sky130_fd_sc_hd__nand2b_1
X_2489_ _3540_/A _2573_/S _2487_/Y _2488_/X vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3211__A1 _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1860_ _1860_/A vssd1 vssd1 vccd1 vccd1 _1860_/Y sky130_fd_sc_hd__inv_2
Xinput12 io_in[26] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
XANTENNA__3202__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 rst_n vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
X_3530_ _3513_/Y _3517_/B _3515_/B vssd1 vssd1 vccd1 vccd1 _3531_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3461_ hold273/X _3470_/B _3460_/Y _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3461_/X sky130_fd_sc_hd__o211a_1
X_3392_ _3635_/A0 hold97/X _3396_/S vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
X_2412_ _2393_/B _2411_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__a21bo_1
X_2343_ _3506_/A _2551_/A _2362_/S vssd1 vssd1 vccd1 vccd1 _2427_/B sky130_fd_sc_hd__mux2_1
X_4013_ _4112_/CLK _4013_/D vssd1 vssd1 vccd1 vccd1 _4013_/Q sky130_fd_sc_hd__dfxtp_1
X_2274_ _1995_/Y _2222_/C _2221_/C _2273_/X vssd1 vssd1 vccd1 vccd1 _2274_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _1989_/A _1996_/S vssd1 vssd1 vccd1 vccd1 _1989_/X sky130_fd_sc_hd__or2_1
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3728_ _3905_/CLK _3728_/D vssd1 vssd1 vccd1 vccd1 _3728_/Q sky130_fd_sc_hd__dfxtp_1
X_3659_ _3507_/A hold316/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1994__A1 _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2943__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output30_A _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2961_ _2967_/A _3824_/Q _3134_/B _3163_/B vssd1 vssd1 vccd1 vccd1 _2961_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1912_ _1906_/A _2180_/B _3506_/A vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__a21o_1
X_2892_ _2962_/A _2992_/A vssd1 vssd1 vccd1 vccd1 _3134_/B sky130_fd_sc_hd__nor2_1
X_1843_ _1843_/A vssd1 vssd1 vccd1 vccd1 _1843_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold615 _4024_/Q vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 _3244_/X vssd1 vssd1 vccd1 vccd1 _3245_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _3297_/X vssd1 vssd1 vccd1 vccd1 _3298_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _3518_/A _3514_/B vssd1 vssd1 vccd1 vccd1 _3513_/Y sky130_fd_sc_hd__nor2_1
X_3444_ _3639_/A0 hold77/X _3444_/S vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__mux2_1
Xhold659 _4017_/Q vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _4020_/Q vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _2992_/Y vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2162__A1 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3375_ _2678_/X _3358_/X _3374_/X vssd1 vssd1 vccd1 vccd1 _3944_/D sky130_fd_sc_hd__a21o_1
X_2326_ _2322_/X _2325_/X _1941_/B _2219_/B vssd1 vssd1 vccd1 vccd1 _2670_/A sky130_fd_sc_hd__a2bb2o_1
X_2257_ _2255_/X _2256_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2261_/C sky130_fd_sc_hd__a21o_1
XANTENNA__3679__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2188_ _2191_/B _2187_/X _2221_/A vssd1 vssd1 vccd1 vccd1 _2189_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout97_A _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2144__A1 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3160_ hold298/X _3165_/B _3159_/Y _3131_/A vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__o211a_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__buf_1
X_3091_ hold623/X _3089_/X _3090_/X _3320_/A vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__a211o_1
X_2111_ _2256_/A _2165_/B _3566_/B vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2042_ _3709_/Q _3721_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3993_ _4014_/CLK _3993_/D vssd1 vssd1 vccd1 vccd1 _3993_/Q sky130_fd_sc_hd__dfxtp_1
X_2944_ _3682_/A0 _2940_/X _2943_/Y vssd1 vssd1 vccd1 vccd1 _2944_/Y sky130_fd_sc_hd__a21oi_1
X_2875_ _2887_/A _2875_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__and3_1
XFILLER_0_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold401 _3899_/Q vssd1 vssd1 vccd1 vccd1 _3261_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _3230_/X vssd1 vssd1 vccd1 vccd1 _3231_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _3760_/Q vssd1 vssd1 vccd1 vccd1 _2789_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _3797_/Q vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _3711_/Q vssd1 vssd1 vccd1 vccd1 _2660_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _3808_/Q vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__clkbuf_4
Xhold456 _3721_/Q vssd1 vssd1 vccd1 vccd1 _2692_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _3783_/Q vssd1 vssd1 vccd1 vccd1 _2843_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3427_ _3604_/C _3455_/A vssd1 vssd1 vccd1 vccd1 _3435_/S sky130_fd_sc_hd__or2_4
Xhold489 _3931_/Q vssd1 vssd1 vccd1 vccd1 _3346_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3640_/A _3358_/B _3640_/C vssd1 vssd1 vccd1 vccd1 _3358_/X sky130_fd_sc_hd__and3_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _1945_/Y _2205_/X _2308_/Y _2616_/A _2181_/Y vssd1 vssd1 vccd1 vccd1 _2309_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3601_/A _3289_/B vssd1 vssd1 vccd1 vccd1 _3911_/D sky130_fd_sc_hd__and2_1
XANTENNA__3399__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2126__A1 _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2660_ _2869_/A _2660_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__and3_1
XFILLER_0_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2591_ _2939_/A _2592_/C vssd1 vssd1 vccd1 vccd1 _2681_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3212_ _1889_/Y _3201_/A _2410_/B _2408_/C vssd1 vssd1 vccd1 vccd1 _3212_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2668__A2 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3143_ _3817_/Q _3199_/B _2971_/X vssd1 vssd1 vccd1 vccd1 _3148_/A sky130_fd_sc_hd__o21ai_4
X_3074_ _2925_/Y _3072_/X _3102_/A _3009_/B _3601_/A vssd1 vssd1 vccd1 vccd1 _3834_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2025_ _3899_/Q _3781_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2025_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3976_ _4073_/CLK _3976_/D vssd1 vssd1 vccd1 vccd1 _3976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2927_ _1925_/C _2925_/Y _2926_/X _3601_/A vssd1 vssd1 vccd1 vccd1 _2927_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1985__B _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2858_ _2658_/X _2853_/X _2857_/X vssd1 vssd1 vccd1 vccd1 _3789_/D sky130_fd_sc_hd__a21o_1
Xhold220 _3623_/X vssd1 vssd1 vccd1 vccd1 _4066_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2789_ _2805_/A _2789_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__and3_1
Xhold231 _3993_/Q vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold253 _3696_/Q vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _2600_/X vssd1 vssd1 vccd1 vccd1 _3700_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _4013_/Q vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _3614_/X vssd1 vssd1 vccd1 vccd1 _4058_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _4098_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _3152_/X vssd1 vssd1 vccd1 vccd1 _3842_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2101__S _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2108__A1 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2659__A2 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2292__B1 _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2044__B1 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2442__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3830_ _4095_/CLK _3830_/D vssd1 vssd1 vccd1 vccd1 _3830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3761_ _3778_/CLK _3761_/D vssd1 vssd1 vccd1 vccd1 _3761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2712_ _3640_/B _2872_/A vssd1 vssd1 vccd1 vccd1 _2741_/S sky130_fd_sc_hd__and2_2
X_3692_ _4011_/CLK _3692_/D vssd1 vssd1 vccd1 vccd1 _3692_/Q sky130_fd_sc_hd__dfxtp_4
X_2643_ _3544_/S _2734_/S _3589_/A _2642_/Y _2640_/B vssd1 vssd1 vccd1 vccd1 _2645_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2574_ _2345_/X _2551_/B _2512_/A vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3126_ _4024_/Q _3124_/Y _3125_/Y _4020_/Q _3097_/Y vssd1 vssd1 vccd1 vccd1 _3126_/X
+ sky130_fd_sc_hd__a221o_1
X_3057_ _3049_/X _3050_/Y _3056_/X _3048_/Y _3022_/X vssd1 vssd1 vccd1 vccd1 _3057_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3471__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2008_ _3600_/B _3658_/A _2008_/C vssd1 vssd1 vccd1 vccd1 _3579_/B sky130_fd_sc_hd__and3b_2
XFILLER_0_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2026__B1 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3959_ _4112_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2290_ _2307_/B _2219_/Y _2287_/X _2205_/X vssd1 vssd1 vccd1 vccd1 _2291_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _4113_/CLK _3813_/D vssd1 vssd1 vccd1 vccd1 _3813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3744_ _4042_/CLK _3744_/D vssd1 vssd1 vccd1 vccd1 _3744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3675_ _3675_/A _3675_/B vssd1 vssd1 vccd1 vccd1 _3683_/S sky130_fd_sc_hd__or2_4
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2626_ _3589_/A _2630_/B hold352/X _2734_/S _1918_/X vssd1 vssd1 vccd1 vccd1 _2626_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3508__B1 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2557_ _3975_/Q _4072_/Q _4064_/Q _4056_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2558_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ hold638/X _2485_/X _3544_/S vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__a21o_1
X_3109_ _3140_/D _3120_/D _3108_/Y _2989_/B vssd1 vssd1 vccd1 vccd1 _3109_/X sky130_fd_sc_hd__a31o_1
X_4089_ _4089_/CLK _4089_/D vssd1 vssd1 vccd1 vccd1 _4089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2722__A1 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 io_in[27] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3460_ _3460_/A _3470_/B vssd1 vssd1 vccd1 vccd1 _3460_/Y sky130_fd_sc_hd__nand2_1
X_2411_ _2406_/X input15/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2411_/X sky130_fd_sc_hd__mux2_1
X_3391_ _3634_/A0 hold11/X _3396_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
X_2342_ _1941_/B _2281_/B _2341_/Y vssd1 vssd1 vccd1 vccd1 _2551_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__2713__B2 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4012_ _4014_/CLK _4012_/D vssd1 vssd1 vccd1 vccd1 _4012_/Q sky130_fd_sc_hd__dfxtp_1
X_2273_ _2192_/A _2192_/B _2192_/C _2194_/A vssd1 vssd1 vccd1 vccd1 _2273_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3727_ _3778_/CLK _3727_/D vssd1 vssd1 vccd1 vccd1 _3727_/Q sky130_fd_sc_hd__dfxtp_1
X_1988_ _1988_/A _2616_/C vssd1 vssd1 vccd1 vccd1 _1988_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2952__A1 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3658_ _3658_/A _3658_/B vssd1 vssd1 vccd1 vccd1 _3674_/S sky130_fd_sc_hd__nand2_8
X_3589_ _3589_/A _3592_/B _3589_/C vssd1 vssd1 vccd1 vccd1 _3589_/Y sky130_fd_sc_hd__nor3_1
X_2609_ _2609_/A _2609_/B vssd1 vssd1 vccd1 vccd1 _2610_/C sky130_fd_sc_hd__or2_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2563__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2943__A1 hold499/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2960_ _2960_/A _3824_/Q _2997_/C vssd1 vssd1 vccd1 vccd1 _3163_/B sky130_fd_sc_hd__and3_2
X_2891_ _2891_/A _2976_/B _3817_/Q _2974_/B vssd1 vssd1 vccd1 vccd1 _3157_/A sky130_fd_sc_hd__or4_4
X_1911_ hold625/X hold269/X _1996_/S vssd1 vssd1 vccd1 vccd1 _3506_/A sky130_fd_sc_hd__mux2_8
X_1842_ _3564_/A vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3512_ hold665/X _3564_/B _3510_/Y _3511_/X _3587_/A vssd1 vssd1 vccd1 vccd1 _3512_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold605 hold739/X vssd1 vssd1 vccd1 vccd1 _3199_/A sky130_fd_sc_hd__clkbuf_2
Xhold627 _3911_/Q vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _3738_/Q vssd1 vssd1 vccd1 vccd1 _2624_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3443_ _1867_/Y hold125/X _3444_/S vssd1 vssd1 vccd1 vccd1 _3443_/X sky130_fd_sc_hd__mux2_1
Xhold638 _3691_/Q vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _2993_/Y vssd1 vssd1 vccd1 vccd1 _3822_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3656_/A _3374_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3374_/X sky130_fd_sc_hd__and3_1
X_2325_ _2289_/Y _2323_/Y _2324_/X _2737_/C vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__o211a_1
X_2256_ _2256_/A _3518_/B vssd1 vssd1 vccd1 vccd1 _2256_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2187_ _3690_/Q _2048_/S _2129_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2187_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2612__B _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2104__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4103_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2536__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _3089_/X _3090_/B _3090_/C vssd1 vssd1 vccd1 vccd1 _3090_/X sky130_fd_sc_hd__and3b_1
X_2110_ _2101_/X _2109_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3566_/B sky130_fd_sc_hd__mux2_2
X_2041_ _2039_/X _2040_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__mux2_1
X_3992_ _4016_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2943_ hold499/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2943_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2874_ _2655_/X _2871_/X _2873_/X vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold402 _3930_/Q vssd1 vssd1 vccd1 vccd1 _3344_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold413 _3750_/Q vssd1 vssd1 vccd1 vccd1 _2767_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 hold732/X vssd1 vssd1 vccd1 vccd1 _2637_/B sky130_fd_sc_hd__clkbuf_2
Xhold424 _3763_/Q vssd1 vssd1 vccd1 vccd1 _2795_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2383__A2 _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold468 _3767_/Q vssd1 vssd1 vccd1 vccd1 _2805_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _3766_/Q vssd1 vssd1 vccd1 vccd1 _2803_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _2693_/X vssd1 vssd1 vccd1 vccd1 _3721_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold479 _3579_/B vssd1 vssd1 vccd1 vccd1 _3564_/B sky130_fd_sc_hd__buf_2
X_3426_ _3874_/Q _3873_/Q vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__nand2b_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _2678_/X _3340_/X _3356_/X vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__a21o_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2308_/A vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__inv_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ input5/X hold627/X _3292_/S vssd1 vssd1 vccd1 vccd1 _3288_/X sky130_fd_sc_hd__mux2_1
X_2239_ _2093_/B _2236_/X _2237_/X _2238_/X vssd1 vssd1 vccd1 vccd1 _2239_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2607__B _3551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2590_ hold559/X _2577_/X _2589_/X _2576_/X _3471_/C1 vssd1 vssd1 vccd1 vccd1 _2590_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3211_ _3691_/Q _3201_/Y _3210_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3211_/X sky130_fd_sc_hd__o211a_1
X_3142_ _3817_/Q _3199_/B _2971_/X vssd1 vssd1 vccd1 vccd1 _3165_/B sky130_fd_sc_hd__o21a_2
XANTENNA__2708__A _3808_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3073_ _3073_/A _3171_/A vssd1 vssd1 vccd1 vccd1 _3102_/A sky130_fd_sc_hd__nor2_1
X_2024_ _2142_/A _2024_/B vssd1 vssd1 vccd1 vccd1 _2024_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ _4072_/CLK _3975_/D vssd1 vssd1 vccd1 vccd1 _3975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3250__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2926_ input4/X _3834_/Q _3072_/B vssd1 vssd1 vccd1 vccd1 _2926_/X sky130_fd_sc_hd__or3_1
XANTENNA__1985__C _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2857_ _2863_/A _2857_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__and3_1
XFILLER_0_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2788_ _2664_/X _2779_/X _2787_/X vssd1 vssd1 vccd1 vccd1 _3759_/D sky130_fd_sc_hd__a21o_1
Xhold210 _3626_/X vssd1 vssd1 vccd1 vccd1 _4069_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _3437_/X vssd1 vssd1 vccd1 vccd1 _3993_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _3946_/Q vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold243 _3949_/Q vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _3465_/X vssd1 vssd1 vccd1 vccd1 _4013_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _2596_/X vssd1 vssd1 vccd1 vccd1 _3696_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _4095_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _3667_/X vssd1 vssd1 vccd1 vccd1 _4098_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold298 _3844_/Q vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _3676_/A0 hold165/X _3416_/S vssd1 vssd1 vccd1 vccd1 _3409_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2513__C1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2044__A1 _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3184__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3760_ _3767_/CLK _3760_/D vssd1 vssd1 vccd1 vccd1 _3760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2711_ _3321_/A _3321_/B _3640_/A vssd1 vssd1 vccd1 vccd1 _2872_/A sky130_fd_sc_hd__and3b_2
X_3691_ _4011_/CLK _3691_/D vssd1 vssd1 vccd1 vccd1 _3691_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2642_ _2642_/A _2642_/B vssd1 vssd1 vccd1 vccd1 _2642_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2573_ _3507_/A _2572_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3299__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2510__A2 _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3125_ _3125_/A _3276_/B vssd1 vssd1 vccd1 vccd1 _3125_/Y sky130_fd_sc_hd__nor2_1
X_3056_ _3055_/X _3056_/B _3056_/C _3056_/D vssd1 vssd1 vccd1 vccd1 _3056_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2007_ _2227_/S _2232_/S vssd1 vssd1 vccd1 vccd1 _2279_/S sky130_fd_sc_hd__or2_2
XANTENNA__2026__A1 _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3958_ _4111_/CLK _3958_/D vssd1 vssd1 vccd1 vccd1 _3958_/Q sky130_fd_sc_hd__dfxtp_1
X_3889_ _4029_/CLK _3889_/D vssd1 vssd1 vccd1 vccd1 _3889_/Q sky130_fd_sc_hd__dfxtp_1
X_2909_ _1841_/Y _3885_/Q _1860_/Y hold665/X vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3526__A1 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout72_A _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2022__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output53_A _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3453__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3812_ _4113_/CLK _3812_/D vssd1 vssd1 vccd1 vccd1 _3812_/Q sky130_fd_sc_hd__dfxtp_1
X_3743_ _3767_/CLK _3743_/D vssd1 vssd1 vccd1 vccd1 _3743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3674_ _2610_/A hold37/X _3674_/S vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__mux2_1
X_2625_ _2732_/A _2732_/B _2624_/A vssd1 vssd1 vccd1 vccd1 _2625_/Y sky130_fd_sc_hd__a21oi_1
X_2556_ _2392_/X _2549_/X _2391_/X vssd1 vssd1 vccd1 vccd1 _2556_/Y sky130_fd_sc_hd__a21oi_1
X_2487_ _2481_/X _2482_/Y _2485_/X _2486_/X vssd1 vssd1 vccd1 vccd1 _2487_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3108_ _3078_/X _3120_/C vssd1 vssd1 vccd1 vccd1 _3108_/Y sky130_fd_sc_hd__nand2b_1
X_4088_ _4088_/CLK _4088_/D vssd1 vssd1 vccd1 vccd1 _4088_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3444__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3039_ _3852_/Q _3043_/A vssd1 vssd1 vccd1 vccd1 _3040_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2107__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3462__A _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3435__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3401__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 io_in[28] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
X_2410_ input1/X _2410_/B _2940_/B vssd1 vssd1 vccd1 vccd1 _2588_/S sky130_fd_sc_hd__and3_4
X_3390_ _3633_/A0 hold169/X _3396_/S vssd1 vssd1 vccd1 vccd1 _3390_/X sky130_fd_sc_hd__mux2_1
X_2341_ _2338_/X _2339_/Y _2340_/X vssd1 vssd1 vccd1 vccd1 _2341_/Y sky130_fd_sc_hd__a21oi_1
X_2272_ _2272_/A _2281_/B vssd1 vssd1 vccd1 vccd1 _2272_/Y sky130_fd_sc_hd__nor2_1
X_4011_ _4011_/CLK _4011_/D vssd1 vssd1 vccd1 vccd1 _4011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ _1987_/A _2180_/B vssd1 vssd1 vccd1 vccd1 _2614_/A sky130_fd_sc_hd__nor2_1
X_3726_ _3905_/CLK _3726_/D vssd1 vssd1 vccd1 vccd1 _3726_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2952__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3657_ _2678_/X _3640_/X _3656_/X vssd1 vssd1 vccd1 vccd1 _4089_/D sky130_fd_sc_hd__a21o_1
X_3588_ _4044_/Q _4043_/Q _2619_/A vssd1 vssd1 vccd1 vccd1 _3589_/C sky130_fd_sc_hd__a21oi_1
X_2608_ _3539_/A _2606_/Y _2607_/X _2573_/S vssd1 vssd1 vccd1 vccd1 _2609_/B sky130_fd_sc_hd__o22a_1
X_2539_ _2564_/A _2538_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2539_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1912__B1 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2563__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3457__A _3467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2943__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2890_ _2891_/A _2976_/B _3817_/Q _2974_/B vssd1 vssd1 vccd1 vccd1 _2890_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__2631__B2 _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1910_ _1987_/A _2616_/C _2158_/S vssd1 vssd1 vccd1 vccd1 _2369_/A sky130_fd_sc_hd__or3_2
XFILLER_0_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1841_ _1841_/A vssd1 vssd1 vccd1 vccd1 _1841_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold606 _2972_/Y vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 hold744/X vssd1 vssd1 vccd1 vccd1 _3050_/A sky130_fd_sc_hd__clkbuf_2
X_3511_ _4044_/Q _3554_/B hold368/X vssd1 vssd1 vccd1 vccd1 _3511_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3442_ _3637_/A0 hold115/X _3444_/S vssd1 vssd1 vccd1 vccd1 _3442_/X sky130_fd_sc_hd__mux2_1
Xhold628 _3288_/X vssd1 vssd1 vccd1 vccd1 _3289_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 _4104_/Q vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _2674_/X _3358_/X _3372_/X vssd1 vssd1 vccd1 vccd1 _3943_/D sky130_fd_sc_hd__a21o_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2235_/Y _2246_/Y _2284_/X _2289_/A _2233_/X vssd1 vssd1 vccd1 vccd1 _2324_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2255_ _2250_/X _2251_/X _2279_/S vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__a21o_1
X_2186_ _3689_/Q _2048_/S _2165_/X _2194_/B vssd1 vssd1 vccd1 vccd1 _2191_/B sky130_fd_sc_hd__a211o_1
Xwrapped_8x305_120 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_120/HI io_out[28] sky130_fd_sc_hd__conb_1
XANTENNA__2870__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3709_ _3795_/CLK _3709_/D vssd1 vssd1 vccd1 vccd1 _3709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3638__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2536__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3629__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2040_ _3929_/Q _3921_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2852__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3991_ _4016_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2942_ _3639_/A0 _2940_/X _2941_/Y vssd1 vssd1 vccd1 vccd1 _2942_/Y sky130_fd_sc_hd__a21oi_1
X_2873_ _2887_/A _2873_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__and3_1
XFILLER_0_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3565__C1 _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3580__A2 _2646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 _3775_/Q vssd1 vssd1 vccd1 vccd1 _2823_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 _3803_/Q vssd1 vssd1 vccd1 vccd1 _2887_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _2796_/X vssd1 vssd1 vccd1 vccd1 _3763_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _3905_/Q vssd1 vssd1 vccd1 vccd1 _3273_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _3800_/Q vssd1 vssd1 vccd1 vccd1 _2881_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 _3749_/Q vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold469 _3724_/Q vssd1 vssd1 vccd1 vccd1 _2698_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3425_ _3639_/A0 hold95/X _3425_/S vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__mux2_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3656_/A _3356_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3356_/X sky130_fd_sc_hd__and3_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2205_/X _2307_/B vssd1 vssd1 vccd1 vccd1 _2308_/A sky130_fd_sc_hd__nand2b_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3601_/A _3287_/B vssd1 vssd1 vccd1 vccd1 _3910_/D sky130_fd_sc_hd__and2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _2238_/A _2238_/B _2238_/C vssd1 vssd1 vccd1 vccd1 _2238_/X sky130_fd_sc_hd__and3_1
X_2169_ _2094_/A _2238_/C _2168_/X _2189_/A vssd1 vssd1 vccd1 vccd1 _2169_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2115__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold499_A _3810_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__A _3695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2598__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2025__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3210_ _1889_/Y _3201_/A _2410_/B _2408_/D vssd1 vssd1 vccd1 vccd1 _3210_/X sky130_fd_sc_hd__a31o_1
X_3141_ hold93/X _3140_/X _3320_/A vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__a21o_1
X_3072_ _3275_/A _3072_/B vssd1 vssd1 vccd1 vccd1 _3072_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2023_ _3710_/Q _3722_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2024_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3974_ _4072_/CLK _3974_/D vssd1 vssd1 vccd1 vccd1 _3974_/Q sky130_fd_sc_hd__dfxtp_1
X_2925_ _3275_/A _3072_/B vssd1 vssd1 vccd1 vccd1 _2925_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2856_ _2655_/X _2853_/X _2855_/X vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 _3976_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
X_2787_ _2805_/A _2787_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2787_/X sky130_fd_sc_hd__and3_1
Xhold200 _3633_/X vssd1 vssd1 vccd1 vccd1 _4075_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _3378_/X vssd1 vssd1 vccd1 vccd1 _3946_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _3381_/X vssd1 vssd1 vccd1 vccd1 _3949_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _4064_/Q vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _4015_/Q vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _3699_/Q vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _3664_/X vssd1 vssd1 vccd1 vccd1 _4095_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _3841_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _3160_/X vssd1 vssd1 vccd1 vccd1 _3844_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3408_ _3874_/Q _3873_/Q _3445_/A vssd1 vssd1 vccd1 vccd1 _3416_/S sky130_fd_sc_hd__or3_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _2678_/X _3322_/X _3338_/X vssd1 vssd1 vccd1 vccd1 _3339_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3404__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2710_ _2834_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _3641_/B sky130_fd_sc_hd__or2_1
X_3690_ _3690_/CLK _3690_/D vssd1 vssd1 vccd1 vccd1 _3690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2641_ _2733_/S _2615_/B _2639_/Y _2640_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _3707_/D
+ sky130_fd_sc_hd__o311a_1
X_2572_ hold559/X _2571_/X _2572_/S vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3124_ _3304_/A _3276_/B vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__nor2_1
X_3055_ _3055_/A _3055_/B _3055_/C _3055_/D vssd1 vssd1 vccd1 vccd1 _3055_/X sky130_fd_sc_hd__or4_1
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2006_ _2227_/S _2573_/S vssd1 vssd1 vccd1 vccd1 _2256_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ _4113_/CLK _3957_/D vssd1 vssd1 vccd1 vccd1 _3957_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3223__A1 _3458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2908_ _4030_/Q _3472_/A _3886_/Q _1840_/Y _2905_/X vssd1 vssd1 vccd1 vccd1 _2918_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3888_ _4092_/CLK _3888_/D vssd1 vssd1 vccd1 vccd1 _3888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ _3269_/A _2839_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout65_A _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3214__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4113_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output46_A _3812_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3811_ _4111_/CLK _3811_/D vssd1 vssd1 vccd1 vccd1 _3811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3742_ _3767_/CLK _3742_/D vssd1 vssd1 vccd1 vccd1 _3742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ _2180_/B hold639/X _3674_/S vssd1 vssd1 vccd1 vccd1 _4104_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2624_ _2624_/A _2624_/B _2732_/B vssd1 vssd1 vccd1 vccd1 _2629_/B sky130_fd_sc_hd__and3_1
XFILLER_0_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2555_ _2392_/A _2553_/X _2554_/X _2612_/B vssd1 vssd1 vccd1 vccd1 _2555_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2486_ _2304_/Y _2430_/B _2508_/A vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3141__B1 _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3107_ _3078_/X _3105_/X _3120_/D _3140_/B vssd1 vssd1 vccd1 vccd1 _3107_/X sky130_fd_sc_hd__a31o_1
X_4087_ _4088_/CLK _4087_/D vssd1 vssd1 vccd1 vccd1 _4087_/Q sky130_fd_sc_hd__dfxtp_1
X_3038_ _4017_/Q _3849_/Q vssd1 vssd1 vccd1 vccd1 _3052_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2123__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3380__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2183__A1 _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 io_in[2] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2033__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2340_ _1945_/Y _2272_/Y _2338_/B _2616_/A _2181_/Y vssd1 vssd1 vccd1 vccd1 _2340_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2271_ _3544_/S _3506_/B _2266_/X _2267_/Y vssd1 vssd1 vccd1 vccd1 _2281_/B sky130_fd_sc_hd__a2bb2o_2
X_4010_ _4016_/CLK _4010_/D vssd1 vssd1 vccd1 vccd1 _4010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1986_ _2610_/A _3596_/A _2393_/B vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__or3_4
XFILLER_0_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3725_ _3902_/CLK _3725_/D vssd1 vssd1 vccd1 vccd1 _3725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3656_ _3656_/A _3656_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3587_ _3587_/A _3587_/B vssd1 vssd1 vccd1 vccd1 _4044_/D sky130_fd_sc_hd__and2_1
X_2607_ _3566_/B _3551_/A _3540_/B _3558_/A vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__or4_1
X_2538_ _4006_/Q _3998_/Q _4014_/Q _3990_/Q _2582_/S1 _3717_/Q vssd1 vssd1 vccd1 vccd1
+ _2538_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2469_ hold9/A hold45/A _4011_/Q hold79/A _2582_/S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1
+ _2469_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2118__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _1840_/A vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__inv_2
X_3510_ _3505_/X _3509_/X _3554_/B vssd1 vssd1 vccd1 vccd1 _3510_/Y sky130_fd_sc_hd__a21oi_1
Xhold618 _3198_/X vssd1 vssd1 vccd1 vccd1 _3861_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold607 _2973_/X vssd1 vssd1 vccd1 vccd1 _3817_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3636_/A0 hold205/X _3444_/S vssd1 vssd1 vccd1 vccd1 _3441_/X sky130_fd_sc_hd__mux2_1
Xhold629 _4046_/Q vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3654_/A _3372_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3372_/X sky130_fd_sc_hd__and3_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2235_/Y _2246_/Y _2284_/X _2233_/X vssd1 vssd1 vccd1 vccd1 _2323_/Y sky130_fd_sc_hd__a31oi_1
X_2254_ _3544_/S _3514_/B vssd1 vssd1 vccd1 vccd1 _2604_/B sky130_fd_sc_hd__or2_2
XANTENNA__3647__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2185_ _2222_/B _2222_/C _2222_/A vssd1 vssd1 vccd1 vccd1 _2189_/B sky130_fd_sc_hd__a21o_1
Xwrapped_8x305_121 vssd1 vssd1 vccd1 vccd1 io_out[2] wrapped_8x305_121/LO sky130_fd_sc_hd__conb_1
XFILLER_0_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1969_ _1988_/A _2180_/B _3554_/A _3540_/A _2616_/B vssd1 vssd1 vccd1 vccd1 _1969_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3708_ _4045_/CLK _3708_/D vssd1 vssd1 vccd1 vccd1 _3708_/Q sky130_fd_sc_hd__dfxtp_1
X_3639_ _3639_/A0 hold39/X _3639_/S vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__mux2_1
XANTENNA__3293__A _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3778_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _4014_/CLK _3990_/D vssd1 vssd1 vccd1 vccd1 _3990_/Q sky130_fd_sc_hd__dfxtp_1
X_2941_ hold512/X _2940_/X _2953_/B1 vssd1 vssd1 vccd1 vccd1 _2941_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2872_ _2872_/A _3358_/B vssd1 vssd1 vccd1 vccd1 _2887_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 _3925_/Q vssd1 vssd1 vccd1 vccd1 _3332_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _3934_/Q vssd1 vssd1 vccd1 vccd1 _3352_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold404 _2888_/X vssd1 vssd1 vccd1 vccd1 _3803_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3424_ _3682_/A0 hold123/X _3425_/S vssd1 vssd1 vccd1 vccd1 _3424_/X sky130_fd_sc_hd__mux2_1
Xhold459 _2882_/X vssd1 vssd1 vccd1 vccd1 _3800_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _2766_/X vssd1 vssd1 vccd1 vccd1 _3749_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _3787_/Q vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3355_ _2674_/X _3340_/X _3354_/X vssd1 vssd1 vccd1 vccd1 _3935_/D sky130_fd_sc_hd__a21o_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2306_/A _2306_/B vssd1 vssd1 vccd1 vccd1 _2313_/A sky130_fd_sc_hd__or2_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3286_ input4/X hold557/X _3292_/S vssd1 vssd1 vccd1 vccd1 _3286_/X sky130_fd_sc_hd__mux2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _2208_/B _2148_/X _1995_/Y vssd1 vssd1 vccd1 vccd1 _2237_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2168_ _2221_/A _2130_/X _2148_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _2168_/X sky130_fd_sc_hd__a31o_1
X_2099_ _3779_/Q _3795_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2099_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2131__S _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout95_A _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2770__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2041__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3140_ _3157_/A _3140_/B _3140_/C _3140_/D vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__or4_1
X_3071_ _3320_/A _3071_/B vssd1 vssd1 vccd1 vccd1 _3833_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2277__A _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2022_ _2020_/X _2021_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3973_ _4073_/CLK _3973_/D vssd1 vssd1 vccd1 vccd1 _3973_/Q sky130_fd_sc_hd__dfxtp_1
X_2924_ _3275_/B _3065_/B _3276_/A _3304_/B vssd1 vssd1 vccd1 vccd1 _3072_/B sky130_fd_sc_hd__or4_4
XFILLER_0_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2855_ _2869_/A _2855_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__and3_1
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2786_ _2661_/X _2779_/X _2785_/X vssd1 vssd1 vccd1 vccd1 _3758_/D sky130_fd_sc_hd__a21o_1
Xhold201 _3703_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _3416_/X vssd1 vssd1 vccd1 vccd1 _3976_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold223 _3975_/Q vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _3620_/X vssd1 vssd1 vccd1 vccd1 _4064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _3469_/X vssd1 vssd1 vccd1 vccd1 _4015_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _2599_/X vssd1 vssd1 vccd1 vccd1 _3699_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _4059_/Q vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _3971_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _3149_/X vssd1 vssd1 vccd1 vccd1 _3841_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _3872_/Q _3871_/Q _3454_/A vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__or3_2
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ _3656_/A _3338_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3338_/X sky130_fd_sc_hd__and3_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3269_/A _3269_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2029__B1 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3465__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2036__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ hold1/X _2640_/B vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__or2_1
X_2571_ _2571_/A _2571_/B _2571_/C _2571_/D vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__and4_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3123_ _3123_/A _3123_/B vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__nand2_1
X_3054_ _3054_/A _3054_/B vssd1 vssd1 vccd1 vccd1 _3055_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ _2238_/A _2005_/B vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__or2_2
XFILLER_0_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3956_ _4111_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
X_2907_ _4039_/Q _1855_/Y _1857_/Y _4034_/Q vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3887_ _4092_/CLK _3887_/D vssd1 vssd1 vccd1 vccd1 _3887_/Q sky130_fd_sc_hd__dfxtp_1
X_2838_ _2655_/X _2835_/Y _2837_/X vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2769_ _2805_/A _2769_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2769_/X sky130_fd_sc_hd__and3_1
XFILLER_0_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2584__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3810_ _4113_/CLK _3810_/D vssd1 vssd1 vccd1 vccd1 _3810_/Q sky130_fd_sc_hd__dfxtp_1
X_3741_ _3791_/CLK _3741_/D vssd1 vssd1 vccd1 vccd1 _3741_/Q sky130_fd_sc_hd__dfxtp_1
X_3672_ _2181_/A _2737_/A _3674_/S vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__mux2_1
X_2623_ _3737_/Q _2726_/B vssd1 vssd1 vccd1 vccd1 _2732_/B sky130_fd_sc_hd__and2_1
X_2554_ _2511_/S _2550_/X _2551_/X _2512_/A vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2716__B2 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2485_ _2483_/X _2570_/B _2570_/A vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__mux2_1
X_3106_ _3106_/A _3118_/B vssd1 vssd1 vccd1 vccd1 _3120_/D sky130_fd_sc_hd__nand2_2
X_4086_ _4088_/CLK _4086_/D vssd1 vssd1 vccd1 vccd1 _4086_/Q sky130_fd_sc_hd__dfxtp_1
X_3037_ _3036_/X _3099_/A _3060_/B vssd1 vssd1 vccd1 vccd1 _3171_/A sky130_fd_sc_hd__and3b_4
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _3939_/CLK _3939_/D vssd1 vssd1 vccd1 vccd1 _3939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2707__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput16 io_in[3] vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__buf_1
XANTENNA__2946__A1 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3371__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2270_ _2266_/B _2266_/C _2269_/X _2646_/B _1867_/Y vssd1 vssd1 vccd1 vccd1 _3506_/B
+ sky130_fd_sc_hd__o32ai_4
XANTENNA__1921__A2 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2557__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1985_ _2616_/B _3540_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2362_/S sky130_fd_sc_hd__and3_4
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3724_ _3795_/CLK _3724_/D vssd1 vssd1 vccd1 vccd1 _3724_/Q sky130_fd_sc_hd__dfxtp_1
X_3655_ _2674_/X _3640_/X _3654_/X vssd1 vssd1 vccd1 vccd1 _4088_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2606_ _2606_/A _2606_/B _2606_/C vssd1 vssd1 vccd1 vccd1 _2606_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_fanout108_A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3586_ _2619_/B _3582_/Y _3585_/X _2613_/Y vssd1 vssd1 vccd1 vccd1 _3587_/B sky130_fd_sc_hd__a22o_1
X_2537_ _2564_/A _2537_/B vssd1 vssd1 vccd1 vccd1 _2537_/Y sky130_fd_sc_hd__nand2b_1
X_2468_ _2585_/A _2468_/B vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1912__A2 _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2399_ _4001_/Q _3993_/Q _4009_/Q hold49/A _2582_/S1 _2582_/S0 vssd1 vssd1 vccd1
+ vccd1 _2399_/X sky130_fd_sc_hd__mux4_1
X_4069_ _4073_/CLK _4069_/D vssd1 vssd1 vccd1 vccd1 _4069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3353__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold608 _3736_/Q vssd1 vssd1 vccd1 vccd1 _2720_/A sky130_fd_sc_hd__buf_1
X_3440_ _3635_/A0 hold113/X _3444_/S vssd1 vssd1 vccd1 vccd1 _3440_/X sky130_fd_sc_hd__mux2_1
Xhold619 hold746/X vssd1 vssd1 vccd1 vccd1 _3584_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3371_ _2671_/X _3358_/X _3370_/X vssd1 vssd1 vccd1 vccd1 _3942_/D sky130_fd_sc_hd__a21o_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _1945_/Y _2288_/B _2289_/A _2616_/A _2181_/Y vssd1 vssd1 vccd1 vccd1 _2322_/X
+ sky130_fd_sc_hd__o221a_1
X_2253_ _2250_/X _2251_/X _2252_/Y _2230_/A _3693_/Q vssd1 vssd1 vccd1 vccd1 _3514_/B
+ sky130_fd_sc_hd__a32o_1
X_2184_ _3692_/Q _2048_/S _2066_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2222_/C sky130_fd_sc_hd__a211o_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1968_ _3321_/A _1948_/X _3321_/B _1967_/X vssd1 vssd1 vccd1 vccd1 _2592_/C sky130_fd_sc_hd__a31oi_4
X_3707_ _4047_/CLK _3707_/D vssd1 vssd1 vccd1 vccd1 _3707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1899_ _1899_/A _1899_/B vssd1 vssd1 vccd1 vccd1 _2610_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3638_ _3682_/A0 hold89/X _3639_/S vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__mux2_1
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3335__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3569_ _2732_/A _3554_/B _3567_/X _3568_/Y hold368/X vssd1 vssd1 vccd1 vccd1 _3569_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2534__C1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2039__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2940_ _2940_/A _2940_/B _3201_/B vssd1 vssd1 vccd1 vccd1 _2940_/X sky130_fd_sc_hd__and3_4
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2871_ _2872_/A _3358_/B vssd1 vssd1 vccd1 vccd1 _2871_/X sky130_fd_sc_hd__and2_2
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2368__A2 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 _3943_/Q vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 _3715_/Q vssd1 vssd1 vccd1 vccd1 _2673_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _3723_/Q vssd1 vssd1 vccd1 vccd1 _2696_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _3927_/Q vssd1 vssd1 vccd1 vccd1 _3336_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _3637_/A0 hold85/X _3425_/S vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__mux2_1
Xhold438 _3765_/Q vssd1 vssd1 vccd1 vccd1 _2801_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3654_/A _3354_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3354_/X sky130_fd_sc_hd__and3_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3830_/Q _3285_/B _3304_/B _3285_/D vssd1 vssd1 vccd1 vccd1 _3292_/S sky130_fd_sc_hd__or4_4
XANTENNA__2738__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2305_ _2349_/B _2369_/B _2303_/X vssd1 vssd1 vccd1 vccd1 _2571_/B sky130_fd_sc_hd__o21a_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2130_/X _2166_/X _2194_/A vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__a21o_1
X_2167_ _2194_/B _2238_/C _2166_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__o211a_1
X_2098_ _3771_/Q _3755_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3253__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2531__A2 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2648__A _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3070_ _3072_/B hold702/X _3058_/X vssd1 vssd1 vccd1 vccd1 _3070_/Y sky130_fd_sc_hd__a21oi_1
X_2021_ _3930_/Q _3922_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3972_ _4081_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2923_ _3123_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _3304_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2854_ _2854_/A _3358_/B vssd1 vssd1 vccd1 vccd1 _2869_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2785_ _2805_/A _2785_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2785_/X sky130_fd_sc_hd__and3_1
Xhold202 _2603_/X vssd1 vssd1 vccd1 vccd1 _3703_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2232__S _2232_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold213 _4109_/Q vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _3415_/X vssd1 vssd1 vccd1 vccd1 _3975_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _4060_/Q vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _3615_/X vssd1 vssd1 vccd1 vccd1 _4059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _4092_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _3411_/X vssd1 vssd1 vccd1 vccd1 _3971_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _3689_/Q vssd1 vssd1 vccd1 vccd1 _3458_/A sky130_fd_sc_hd__buf_2
X_3406_ _3639_/A0 hold173/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3406_/X sky130_fd_sc_hd__mux2_1
X_3337_ _2674_/X _3322_/X _3336_/X vssd1 vssd1 vccd1 vccd1 _3927_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3571__B _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _2667_/X _3257_/Y _3267_/X vssd1 vssd1 vccd1 vccd1 _3902_/D sky130_fd_sc_hd__a21o_1
X_2219_ _3652_/B _2219_/B vssd1 vssd1 vccd1 vccd1 _2219_/Y sky130_fd_sc_hd__nand2b_1
X_3199_ _3199_/A _3199_/B vssd1 vssd1 vccd1 vccd1 _3199_/X sky130_fd_sc_hd__and2_1
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2052__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2570_ _2570_/A _2570_/B vssd1 vssd1 vccd1 vccd1 _2572_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3122_ _3157_/A _2988_/B _3307_/C _3117_/X _3116_/X vssd1 vssd1 vccd1 vccd1 _3130_/S
+ sky130_fd_sc_hd__o311a_1
X_3053_ _3053_/A _3053_/B _3053_/C _3053_/D vssd1 vssd1 vccd1 vccd1 _3055_/C sky130_fd_sc_hd__or4_1
X_2004_ _2238_/A _2005_/B vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3955_ _4112_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2906_ _1844_/Y _3882_/Q _1859_/Y _4032_/Q vssd1 vssd1 vccd1 vccd1 _2906_/X sky130_fd_sc_hd__a22o_1
X_3886_ _4092_/CLK _3886_/D vssd1 vssd1 vccd1 vccd1 _3886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2837_ _3269_/A _2837_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__and3_1
X_2768_ _2661_/X _2761_/X _2767_/X vssd1 vssd1 vccd1 vccd1 _3750_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2699_ _2664_/X _2690_/Y _2698_/X vssd1 vssd1 vccd1 vccd1 _3724_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_13_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3447__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3521__S _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2926__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2137__S _2155_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2489__A1 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2584__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3438__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ _3803_/CLK _3740_/D vssd1 vssd1 vccd1 vccd1 _3740_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3610__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3671_ _3554_/A hold328/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3671_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _4047_/Q _4046_/Q _3736_/Q _3592_/B vssd1 vssd1 vccd1 vccd1 _2726_/B sky130_fd_sc_hd__and4_1
X_2553_ _3506_/A _2573_/S _2550_/X _2552_/X vssd1 vssd1 vccd1 vccd1 _2553_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1915__A _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2484_ _2484_/A _2484_/B vssd1 vssd1 vccd1 vccd1 _2570_/B sky130_fd_sc_hd__or2_1
XANTENNA__3677__A0 _1862_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3429__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4085_ _4088_/CLK _4085_/D vssd1 vssd1 vccd1 vccd1 _4085_/Q sky130_fd_sc_hd__dfxtp_1
X_3105_ _3134_/C _3140_/D vssd1 vssd1 vccd1 vccd1 _3105_/X sky130_fd_sc_hd__or2_1
X_3036_ _3833_/Q _3036_/B _3099_/C vssd1 vssd1 vccd1 vccd1 _3036_/X sky130_fd_sc_hd__or3_1
XFILLER_0_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3938_ _3938_/CLK _3938_/D vssd1 vssd1 vccd1 vccd1 _3938_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2955__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3869_ _4014_/CLK _3869_/D vssd1 vssd1 vccd1 vccd1 _3869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3938_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3668__A0 _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2643__A1 _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2396__C_N input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 io_in[4] vssd1 vssd1 vccd1 vccd1 _1886_/A sky130_fd_sc_hd__buf_1
XANTENNA__2946__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3659__A0 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2557__S1 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output51_A _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2882__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1984_ _2008_/C _3600_/B vssd1 vssd1 vccd1 vccd1 _2393_/B sky130_fd_sc_hd__nand2b_4
XFILLER_0_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3723_ _3795_/CLK _3723_/D vssd1 vssd1 vccd1 vccd1 _3723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3654_ _3654_/A _3654_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2605_ _3502_/B _3525_/B _3518_/B _2277_/X _2604_/X vssd1 vssd1 vccd1 vccd1 _2609_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3585_ _2619_/B _3584_/Y _3589_/A _3506_/A vssd1 vssd1 vccd1 vccd1 _3585_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2536_ _3974_/Q _4071_/Q _4063_/Q hold23/A _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2537_/B sky130_fd_sc_hd__mux4_1
X_2467_ _3971_/Q _4068_/Q _4060_/Q _4052_/Q _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2468_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2398_ _2564_/A _2398_/B vssd1 vssd1 vccd1 vccd1 _2398_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _4073_/CLK _4068_/D vssd1 vssd1 vccd1 vccd1 _4068_/Q sky130_fd_sc_hd__dfxtp_1
X_3019_ _3050_/C _3019_/B vssd1 vssd1 vccd1 vccd1 _3048_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2864__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold609 _3692_/Q vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3370_ _3654_/A _3370_/B _3374_/C vssd1 vssd1 vccd1 vccd1 _3370_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2060__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _2571_/C vssd1 vssd1 vccd1 vccd1 _2508_/A sky130_fd_sc_hd__inv_2
X_2252_ _2424_/A _2424_/B _2230_/A vssd1 vssd1 vccd1 vccd1 _2252_/Y sky130_fd_sc_hd__a21oi_1
X_2183_ _3691_/Q _2048_/S _2147_/X _2194_/B vssd1 vssd1 vccd1 vccd1 _2222_/B sky130_fd_sc_hd__a211o_1
XANTENNA__2296__A _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3568__C1 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ _4047_/CLK _3706_/D vssd1 vssd1 vccd1 vccd1 _3706_/Q sky130_fd_sc_hd__dfxtp_1
X_1967_ _3913_/Q _1929_/Y _3321_/B _1957_/Y _1966_/X vssd1 vssd1 vccd1 vccd1 _1967_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1898_ _1899_/A _1899_/B vssd1 vssd1 vccd1 vccd1 _2616_/B sky130_fd_sc_hd__or2_2
X_3637_ _3637_/A0 hold135/X _3639_/S vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3568_ _3559_/B _3562_/X _3566_/Y _1988_/Y _3554_/A vssd1 vssd1 vccd1 vccd1 _3568_/Y
+ sky130_fd_sc_hd__a311oi_1
X_2519_ _3981_/Q _4110_/Q _3965_/Q _3957_/Q _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2520_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_11_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3499_ _3554_/B _3499_/B vssd1 vssd1 vccd1 vccd1 _3499_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2846__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3574__A2 _2646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4092_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3262__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2055__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2870_ _2678_/X _2853_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold406 _3801_/Q vssd1 vssd1 vccd1 vccd1 _2883_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _3770_/Q vssd1 vssd1 vccd1 vccd1 _2811_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3422_ _3636_/A0 hold141/X _3425_/S vssd1 vssd1 vccd1 vccd1 _3422_/X sky130_fd_sc_hd__mux2_1
Xhold428 _3935_/Q vssd1 vssd1 vccd1 vccd1 _3354_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold439 _2802_/X vssd1 vssd1 vccd1 vccd1 _3765_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _2671_/X _3340_/X _3352_/X vssd1 vssd1 vccd1 vccd1 _3934_/D sky130_fd_sc_hd__a21o_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3284_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3909_/D sky130_fd_sc_hd__and2_1
X_2304_ _2349_/B _2369_/B _2303_/X vssd1 vssd1 vccd1 vccd1 _2304_/Y sky130_fd_sc_hd__o21ai_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _2285_/A vssd1 vssd1 vccd1 vccd1 _2235_/Y sky130_fd_sc_hd__inv_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2166_ _3689_/Q _2048_/S _2165_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2166_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2754__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2097_ _2095_/X _2096_/X _2151_/S vssd1 vssd1 vccd1 vccd1 _2097_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2999_ _3199_/B _3163_/B _2997_/Y _2967_/A _3320_/A vssd1 vssd1 vccd1 vccd1 _2999_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold547_A _3813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2452__C1 _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2020_ _4083_/Q _3938_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__mux2_1
X_3971_ _4072_/CLK _3971_/D vssd1 vssd1 vccd1 vccd1 _3971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2922_ _3065_/B _3276_/A vssd1 vssd1 vccd1 vccd1 _2922_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2853_ _2854_/A _3358_/B vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__and2_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2784_ _2658_/X _2779_/X _2783_/X vssd1 vssd1 vccd1 vccd1 _2784_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold214 _3679_/X vssd1 vssd1 vccd1 vccd1 _4109_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _4006_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _4056_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _4091_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _3661_/X vssd1 vssd1 vccd1 vccd1 _4092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _3891_/Q vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _3616_/X vssd1 vssd1 vccd1 vccd1 _4060_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ _3682_/A0 hold143/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3405_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3336_ _3654_/A _3336_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3336_/X sky130_fd_sc_hd__and3_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3269_/A _3267_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3267_/X sky130_fd_sc_hd__and3_1
X_2218_ _4087_/Q _2219_/B vssd1 vssd1 vccd1 vccd1 _2288_/A sky130_fd_sc_hd__and2b_1
X_3198_ _3050_/A _3189_/S _3197_/X _3497_/A vssd1 vssd1 vccd1 vccd1 _3198_/X sky130_fd_sc_hd__o211a_1
X_2149_ hold7/A _3802_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3121_ _3120_/Y _3121_/B _3308_/A vssd1 vssd1 vccd1 vccd1 _3307_/C sky130_fd_sc_hd__nand3b_1
X_3052_ hold3/A _3052_/B _3052_/C _3171_/A vssd1 vssd1 vccd1 vccd1 _3053_/D sky130_fd_sc_hd__or4b_1
XANTENNA__3456__A1 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2003_ _2194_/A _2192_/A vssd1 vssd1 vccd1 vccd1 _2005_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3208__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3954_ _4113_/CLK _3954_/D vssd1 vssd1 vccd1 vccd1 _3954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3885_ _4031_/CLK _3885_/D vssd1 vssd1 vccd1 vccd1 _3885_/Q sky130_fd_sc_hd__dfxtp_1
X_2905_ _4042_/Q _1852_/Y _1858_/Y _4033_/Q vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__a22o_1
X_2836_ _3258_/A _3359_/B vssd1 vssd1 vccd1 vccd1 _2851_/C sky130_fd_sc_hd__or2_2
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3392__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2767_ _2805_/A _2767_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2767_/X sky130_fd_sc_hd__and3_1
X_2698_ _2698_/A _2698_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__and3_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ hold718/X _3314_/S _3308_/Y _3318_/X vssd1 vssd1 vccd1 vccd1 _3319_/X sky130_fd_sc_hd__o22a_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2153__S _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3383__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2949__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _1959_/D hold563/X _3674_/S vssd1 vssd1 vccd1 vccd1 _3670_/X sky130_fd_sc_hd__mux2_1
X_2621_ _2621_/A _3592_/A _3592_/B vssd1 vssd1 vccd1 vccd1 _2720_/B sky130_fd_sc_hd__nand3_1
X_2552_ hold520/X _2549_/X _1930_/Y vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2483_ _2369_/A _2369_/B _2420_/Y _2424_/X vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__a31o_1
X_3104_ _3828_/Q _3118_/B _3120_/A vssd1 vssd1 vccd1 vccd1 _3140_/D sky130_fd_sc_hd__or3b_1
X_4084_ _4089_/CLK _4084_/D vssd1 vssd1 vccd1 vccd1 _4084_/Q sky130_fd_sc_hd__dfxtp_1
X_3035_ _3853_/Q _3040_/A vssd1 vssd1 vccd1 vccd1 _3041_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2762__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3577__B _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3937_ _3939_/CLK _3937_/D vssd1 vssd1 vccd1 vccd1 _3937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3868_ _4103_/CLK _3868_/D vssd1 vssd1 vccd1 vccd1 _3868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3799_ _4042_/CLK _3799_/D vssd1 vssd1 vccd1 vccd1 _3799_/Q sky130_fd_sc_hd__dfxtp_1
X_2819_ _2863_/A _2819_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2819_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3532__S _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2340__B2 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2340__A1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 io_in[5] vssd1 vssd1 vccd1 vccd1 _1885_/A sky130_fd_sc_hd__buf_1
XANTENNA__2331__A1 _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output44_A _3810_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1983_ _2008_/C _3600_/B vssd1 vssd1 vccd1 vccd1 _2612_/B sky130_fd_sc_hd__and2b_4
X_3722_ _3902_/CLK _3722_/D vssd1 vssd1 vccd1 vccd1 _3722_/Q sky130_fd_sc_hd__dfxtp_1
X_3653_ _2671_/X _3640_/X _3652_/X vssd1 vssd1 vccd1 vccd1 _4087_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_70_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2604_ _3529_/B _2604_/B _3506_/B _3507_/B vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__or4_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3584_ _3584_/A _3596_/B vssd1 vssd1 vccd1 vccd1 _3584_/Y sky130_fd_sc_hd__nand2_1
X_2535_ _2393_/X _2529_/B _2390_/Y vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2466_ _2393_/X _2458_/X _2390_/Y vssd1 vssd1 vccd1 vccd1 _2466_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2322__B2 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2322__A1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2397_ _3969_/Q _4066_/Q _4058_/Q _4050_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2398_/B sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4067_ _4072_/CLK _4067_/D vssd1 vssd1 vccd1 vccd1 _4067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3018_ _3193_/A _3024_/B _3195_/A vssd1 vssd1 vccd1 vccd1 _3019_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3498__A _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _3321_/A _2319_/X _2362_/S vssd1 vssd1 vccd1 vccd1 _2571_/C sky130_fd_sc_hd__mux2_2
X_2251_ _2220_/A _2195_/X _2191_/X _2093_/B vssd1 vssd1 vccd1 vccd1 _2251_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2296__B _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2182_ _1945_/Y _2177_/Y _2291_/A _2616_/A _2181_/Y vssd1 vssd1 vccd1 vccd1 _2182_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4080_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1966_ _3602_/A _4098_/Q _2647_/A vssd1 vssd1 vccd1 vccd1 _1966_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _4045_/CLK _3705_/D vssd1 vssd1 vccd1 vccd1 _3705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1897_ _3602_/A _3600_/B _3909_/Q vssd1 vssd1 vccd1 vccd1 _1899_/B sky130_fd_sc_hd__nor3_2
XANTENNA_fanout113_A input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3636_ _3636_/A0 hold117/X _3639_/S vssd1 vssd1 vccd1 vccd1 _3636_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3567_ _3559_/B _3562_/X _3566_/Y vssd1 vssd1 vccd1 vccd1 _3567_/X sky130_fd_sc_hd__a21o_1
X_2518_ _2585_/A _2517_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3498_ _3507_/A _3498_/B vssd1 vssd1 vccd1 vccd1 _3499_/B sky130_fd_sc_hd__xnor2_1
X_2449_ _1886_/Y _2448_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2782__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2161__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2071__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 _3741_/Q vssd1 vssd1 vccd1 vccd1 _2746_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _3727_/Q vssd1 vssd1 vccd1 vccd1 _2704_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _3635_/A0 hold41/X _3425_/S vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
Xhold429 _3791_/Q vssd1 vssd1 vccd1 vccd1 _2861_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3352_ _3352_/A _3352_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3352_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2303_ _2834_/A _2362_/S vssd1 vssd1 vccd1 vccd1 _2303_/X sky130_fd_sc_hd__or2_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ input7/X hold661/X _3283_/S vssd1 vssd1 vccd1 vccd1 _3283_/X sky130_fd_sc_hd__mux2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _4086_/Q _2234_/B vssd1 vssd1 vccd1 vccd1 _2285_/A sky130_fd_sc_hd__xnor2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _2256_/A _2165_/B _3558_/A vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__and3_1
X_2096_ _3747_/Q _3763_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2096_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2998_ _3131_/A _2998_/B _2998_/C vssd1 vssd1 vccd1 vccd1 _2998_/X sky130_fd_sc_hd__and3_1
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1949_ _1949_/A _1996_/S vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__or2_2
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2764__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3619_ _1866_/Y hold149/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3619_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2010__A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2156__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2755__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _4081_/CLK _3970_/D vssd1 vssd1 vccd1 vccd1 _3970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2921_ _3100_/A _3060_/B vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2852_ _2678_/X _2835_/Y _2851_/X vssd1 vssd1 vccd1 vccd1 _3787_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2783_ _2805_/A _2783_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__and3_1
Xhold215 _3990_/Q vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _3451_/X vssd1 vssd1 vccd1 vccd1 _4006_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _3611_/X vssd1 vssd1 vccd1 vccd1 _4056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 _4062_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _3250_/X vssd1 vssd1 vccd1 vccd1 _3891_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold237 _3973_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _3637_/A0 hold197/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3404_/X sky130_fd_sc_hd__mux2_1
X_3335_ _2671_/X _3322_/X _3334_/X vssd1 vssd1 vccd1 vccd1 _3926_/D sky130_fd_sc_hd__a21o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _2664_/X _3257_/Y _3265_/X vssd1 vssd1 vccd1 vccd1 _3901_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3459__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _3544_/S _2606_/C _2213_/X vssd1 vssd1 vccd1 vccd1 _2219_/B sky130_fd_sc_hd__o21a_1
X_3197_ _3861_/Q _3197_/B vssd1 vssd1 vccd1 vccd1 _3197_/X sky130_fd_sc_hd__or2_1
X_2148_ _3691_/Q _2048_/S _2147_/X _2192_/A vssd1 vssd1 vccd1 vccd1 _2148_/X sky130_fd_sc_hd__a211o_1
X_2079_ _2142_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _2079_/X sky130_fd_sc_hd__or2_1
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3120_ _3120_/A _3140_/B _3120_/C _3120_/D vssd1 vssd1 vccd1 vccd1 _3120_/Y sky130_fd_sc_hd__nor4_1
X_3051_ _4021_/Q _3051_/B vssd1 vssd1 vccd1 vccd1 _3053_/C sky130_fd_sc_hd__xnor2_1
X_2002_ _2194_/A _2192_/A vssd1 vssd1 vccd1 vccd1 _2220_/A sky130_fd_sc_hd__nand2_1
XANTENNA__1920__C _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3953_ _4111_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
X_2904_ _3099_/C _3304_/A vssd1 vssd1 vccd1 vccd1 _2937_/A sky130_fd_sc_hd__or2_1
X_3884_ _4092_/CLK _3884_/D vssd1 vssd1 vccd1 vccd1 _3884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2835_ _3258_/A _3359_/B vssd1 vssd1 vccd1 vccd1 _2835_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__2719__B2 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2766_ _2658_/X _2761_/X _2765_/X vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__a21o_1
X_2697_ _2661_/X _2690_/Y _2696_/X vssd1 vssd1 vccd1 vccd1 _3723_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2578__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3316_/X _3317_/X _2988_/B vssd1 vssd1 vccd1 vccd1 _3318_/X sky130_fd_sc_hd__o21a_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3676_/A0 hold73/X _3256_/S vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__mux2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold590 _3855_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2620_ _3592_/A _3592_/B vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2551_ _2551_/A _2551_/B vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__and2_1
X_2482_ _2304_/Y _2427_/X _2428_/X _2508_/A vssd1 vssd1 vccd1 vccd1 _2482_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__2334__C1 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4083_ _4088_/CLK _4083_/D vssd1 vssd1 vccd1 vccd1 _4083_/Q sky130_fd_sc_hd__dfxtp_2
X_3103_ _3169_/B _3057_/X _3102_/X _2988_/B _3199_/B vssd1 vssd1 vccd1 vccd1 _3103_/X
+ sky130_fd_sc_hd__o311a_1
X_3034_ _4022_/Q _3854_/Q vssd1 vssd1 vccd1 vccd1 _3054_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3936_ _3939_/CLK _3936_/D vssd1 vssd1 vccd1 vccd1 _3936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3867_ _4072_/CLK _3867_/D vssd1 vssd1 vccd1 vccd1 _3867_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ _4042_/CLK _3798_/D vssd1 vssd1 vccd1 vccd1 _3798_/Q sky130_fd_sc_hd__dfxtp_1
X_2818_ _2655_/X _2815_/X _2817_/X vssd1 vssd1 vccd1 vccd1 _2818_/X sky130_fd_sc_hd__a21o_1
X_2749_ _2661_/X _2742_/X _2748_/X vssd1 vssd1 vccd1 vccd1 _3742_/D sky130_fd_sc_hd__a21o_1
XANTENNA__3365__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2325__C1 _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3791_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 io_in[6] vssd1 vssd1 vccd1 vccd1 _1884_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3292__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2074__S _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1982_ _3554_/A _2268_/A vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3721_ _3795_/CLK _3721_/D vssd1 vssd1 vccd1 vccd1 _3721_/Q sky130_fd_sc_hd__dfxtp_1
X_3652_ _3654_/A _3652_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__and3_1
XANTENNA__3347__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3583_ _3584_/A _2613_/Y _3581_/Y _3582_/Y _3587_/A vssd1 vssd1 vccd1 vccd1 _4043_/D
+ sky130_fd_sc_hd__o221a_1
X_2603_ _3639_/A0 hold201/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2555__C1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2534_ _2392_/A _2531_/X _2533_/X _2612_/B vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2465_ _2511_/S _2460_/X _2464_/Y _2512_/A vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2396_ _2592_/C _2592_/B input2/X vssd1 vssd1 vccd1 vccd1 _2587_/S sky130_fd_sc_hd__nor3b_4
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4066_ _4073_/CLK _4066_/D vssd1 vssd1 vccd1 vccd1 _4066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3017_ _3195_/A _3193_/A _3024_/B vssd1 vssd1 vccd1 vccd1 _3050_/C sky130_fd_sc_hd__and3_1
XANTENNA__3283__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3919_ _4080_/CLK _3919_/D vssd1 vssd1 vccd1 vccd1 _3919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2159__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1998__S _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3329__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _2248_/X _2249_/X _2238_/B vssd1 vssd1 vccd1 vccd1 _2250_/X sky130_fd_sc_hd__a21o_1
X_2181_ _2181_/A _2616_/C vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__nand2_2
Xwrapped_8x305_114 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_114/HI io_out[22] sky130_fd_sc_hd__conb_1
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1965_ _2410_/B vssd1 vssd1 vccd1 vccd1 _2939_/B sky130_fd_sc_hd__inv_2
X_3704_ _4042_/CLK _3704_/D vssd1 vssd1 vccd1 vccd1 _3704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1896_ _3602_/A _3600_/B hold37/X vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__o21ba_2
X_3635_ _3635_/A0 hold57/X _3639_/S vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout106_A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3566_ _3566_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _3566_/Y sky130_fd_sc_hd__xnor2_1
X_2517_ _4005_/Q _3997_/Q _4013_/Q hold53/A _2582_/S1 _2582_/S0 vssd1 vssd1 vccd1
+ vccd1 _2517_/X sky130_fd_sc_hd__mux4_1
X_3497_ _3497_/A _3497_/B vssd1 vssd1 vccd1 vccd1 _4029_/D sky130_fd_sc_hd__and2_1
X_2448_ _3720_/Q _2445_/Y _2447_/Y _2441_/Y _2443_/Y vssd1 vssd1 vccd1 vccd1 _2448_/X
+ sky130_fd_sc_hd__a32o_1
X_2379_ _2378_/X _2377_/Y _2484_/A vssd1 vssd1 vccd1 vccd1 _2507_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3256__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4049_ _4105_/CLK _4049_/D vssd1 vssd1 vccd1 vccd1 _4049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2231__A1 _3691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold408 _2747_/X vssd1 vssd1 vccd1 vccd1 _3741_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _3634_/A0 hold91/X _3425_/S vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__mux2_1
Xhold419 _3938_/Q vssd1 vssd1 vccd1 vccd1 _3362_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3351_ _2667_/X _3340_/X _3350_/X vssd1 vssd1 vccd1 vccd1 _3933_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2302_ _2834_/A _2296_/X _2297_/X _2194_/A vssd1 vssd1 vccd1 vccd1 _2369_/B sky130_fd_sc_hd__o22a_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3601_/A _3282_/B vssd1 vssd1 vccd1 vccd1 _3908_/D sky130_fd_sc_hd__and2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _4086_/Q _2234_/B vssd1 vssd1 vccd1 vccd1 _2233_/X sky130_fd_sc_hd__and2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2164_ _2155_/X _2163_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3558_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2095_ hold35/A _3803_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2095_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2461__A1 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2997_ _2997_/A _3199_/B _2997_/C vssd1 vssd1 vccd1 vccd1 _2997_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3410__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1948_ _3322_/A _2296_/B _1948_/C vssd1 vssd1 vccd1 vccd1 _1948_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1879_ _3656_/B vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ _3636_/A0 hold259/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3618_/X sky130_fd_sc_hd__mux2_1
X_3549_ _3540_/A _3540_/B _3548_/X vssd1 vssd1 vccd1 vccd1 _3553_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2452__A1 _3458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3401__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2204__A1 _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2920_ _2910_/X hold716/X _2919_/Y _3275_/C vssd1 vssd1 vccd1 vccd1 _3065_/B sky130_fd_sc_hd__a31o_2
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2851_ _3656_/A _2851_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2851_/X sky130_fd_sc_hd__and3_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2782_ _2655_/X _2779_/X _2781_/X vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold205 _3997_/Q vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 _3433_/X vssd1 vssd1 vccd1 vccd1 _3990_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3403_ _3636_/A0 hold229/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3403_/X sky130_fd_sc_hd__mux2_1
Xhold249 _4038_/Q vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__buf_1
Xhold227 _3948_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _3413_/X vssd1 vssd1 vccd1 vccd1 _3973_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3334_ _3654_/A _3334_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3334_/X sky130_fd_sc_hd__and3_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3269_/A _3265_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3265_/X sky130_fd_sc_hd__and3_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _3634_/A0 _2646_/B _2211_/Y _2215_/X vssd1 vssd1 vccd1 vccd1 _2606_/C sky130_fd_sc_hd__o22a_1
X_3196_ _4028_/Q _3189_/S _3195_/X _3114_/A vssd1 vssd1 vccd1 vccd1 _3196_/X sky130_fd_sc_hd__o211a_1
X_2147_ _2256_/A _2165_/B _3540_/B vssd1 vssd1 vccd1 vccd1 _2147_/X sky130_fd_sc_hd__and3_1
X_2078_ _3711_/Q _3723_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2079_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2781__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3050_ _3050_/A _3861_/Q _3050_/C vssd1 vssd1 vccd1 vccd1 _3050_/Y sky130_fd_sc_hd__nor3_1
X_2001_ _2194_/A _2192_/A vssd1 vssd1 vccd1 vccd1 _2238_/A sky130_fd_sc_hd__and2_1
XANTENNA__2077__S _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3952_ _4080_/CLK _3952_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3883_ _4031_/CLK _3883_/D vssd1 vssd1 vccd1 vccd1 _3883_/Q sky130_fd_sc_hd__dfxtp_1
X_2903_ _3099_/C _3304_/A vssd1 vssd1 vccd1 vccd1 _3169_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2106__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2834_ _2834_/A _2834_/B vssd1 vssd1 vccd1 vccd1 _3359_/B sky130_fd_sc_hd__or2_1
XFILLER_0_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1945__A _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2765_ _2805_/A _2765_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__and3_1
XFILLER_0_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2696_ _2698_/A _2696_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__and3_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2578__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ hold597/X _3124_/Y _3304_/Y hold571/X vssd1 vssd1 vccd1 vccd1 _3317_/X sky130_fd_sc_hd__a22o_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3631_/A _3872_/Q _3871_/Q vssd1 vssd1 vccd1 vccd1 _3256_/S sky130_fd_sc_hd__or3b_4
X_3179_ _3179_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3179_/X sky130_fd_sc_hd__or2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2450__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold580 _4096_/Q vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2343__A0 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 _3185_/X vssd1 vssd1 vccd1 vccd1 _3186_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2949__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2550_ _2549_/X _2550_/B _2571_/C _2571_/B vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__and4b_1
X_2481_ _2571_/A _2333_/Y _2416_/Y _2304_/Y vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3102_ _3102_/A _3102_/B _3115_/B _3102_/D vssd1 vssd1 vccd1 vccd1 _3102_/X sky130_fd_sc_hd__and4_1
X_4082_ _4089_/CLK _4082_/D vssd1 vssd1 vccd1 vccd1 _4082_/Q sky130_fd_sc_hd__dfxtp_1
X_3033_ _4023_/Q _3033_/B vssd1 vssd1 vccd1 vccd1 _3055_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2496__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ _3938_/CLK _3935_/D vssd1 vssd1 vccd1 vccd1 _3935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3866_ _4072_/CLK _3866_/D vssd1 vssd1 vccd1 vccd1 _3866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ _4045_/CLK _3797_/D vssd1 vssd1 vccd1 vccd1 _3797_/Q sky130_fd_sc_hd__dfxtp_1
X_2817_ _2869_/A _2817_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__and3_1
X_2748_ _2805_/A _2748_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__and3_1
XANTENNA__2573__A0 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2679_ _2652_/Y _2678_/X _2676_/X vssd1 vssd1 vccd1 vccd1 _3716_/D sky130_fd_sc_hd__a21o_1
XANTENNA__2876__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2800__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1981_ hold589/X _1890_/Y _1979_/X vssd1 vssd1 vccd1 vccd1 _2378_/A sky130_fd_sc_hd__o21a_2
X_3720_ _4014_/CLK _3720_/D vssd1 vssd1 vccd1 vccd1 _3720_/Q sky130_fd_sc_hd__dfxtp_4
X_3651_ _2667_/X _3640_/X _3650_/X vssd1 vssd1 vccd1 vccd1 _4086_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3582_ _3584_/A _3589_/A _2613_/Y vssd1 vssd1 vccd1 vccd1 _3582_/Y sky130_fd_sc_hd__o21ai_1
X_2602_ _3682_/A0 hold181/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__mux2_1
X_2533_ _2511_/S _2529_/X _2532_/X vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2464_ _2670_/A _2511_/S vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2858__A1 _2658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2395_ _3878_/Q _3877_/Q _3876_/Q _3875_/Q vssd1 vssd1 vccd1 vccd1 _2592_/B sky130_fd_sc_hd__or4_2
X_4065_ _4073_/CLK _4065_/D vssd1 vssd1 vccd1 vccd1 _4065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3016_ _3858_/Q _3027_/A vssd1 vssd1 vccd1 vccd1 _3024_/B sky130_fd_sc_hd__and2_1
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2469__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3918_ _4095_/CLK _3918_/D vssd1 vssd1 vccd1 vccd1 _3918_/Q sky130_fd_sc_hd__dfxtp_1
X_3849_ _4029_/CLK _3849_/D vssd1 vssd1 vccd1 vccd1 _3849_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3274__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _2616_/A _2180_/B vssd1 vssd1 vccd1 vccd1 _2737_/C sky130_fd_sc_hd__nor2_2
Xwrapped_8x305_115 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_115/HI io_out[23] sky130_fd_sc_hd__conb_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1964_ _3321_/A _1948_/X _1954_/Y _1963_/X vssd1 vssd1 vccd1 vccd1 _2410_/B sky130_fd_sc_hd__a31o_4
X_3703_ _4080_/CLK _3703_/D vssd1 vssd1 vccd1 vccd1 _3703_/Q sky130_fd_sc_hd__dfxtp_1
X_3634_ _3634_/A0 hold139/X _3639_/S vssd1 vssd1 vccd1 vccd1 _3634_/X sky130_fd_sc_hd__mux2_1
X_1895_ _1895_/A _1895_/B vssd1 vssd1 vccd1 vccd1 _2181_/A sky130_fd_sc_hd__and2_2
X_3565_ hold368/X _3563_/X _3564_/X _3658_/B vssd1 vssd1 vccd1 vccd1 _4036_/D sky130_fd_sc_hd__o211a_1
X_3496_ hold652/X _3050_/A _3496_/S vssd1 vssd1 vccd1 vccd1 _3497_/B sky130_fd_sc_hd__mux2_1
X_2516_ _2564_/A _2516_/B vssd1 vssd1 vccd1 vccd1 _2516_/Y sky130_fd_sc_hd__nand2b_1
X_2447_ _2585_/A _2447_/B vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2378_ _2378_/A _2378_/B _2378_/C vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__or3_1
X_4048_ _4105_/CLK _4048_/D vssd1 vssd1 vccd1 vccd1 _4048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2024__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1863__A _3460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 _3939_/Q vssd1 vssd1 vccd1 vccd1 _3364_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3350_ _3352_/A _3350_/B _3356_/C vssd1 vssd1 vccd1 vccd1 _3350_/X sky130_fd_sc_hd__and3_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _3566_/A _2349_/B vssd1 vssd1 vccd1 vccd1 _2301_/Y sky130_fd_sc_hd__nand2_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3281_ input6/X _1902_/C _3283_/S vssd1 vssd1 vccd1 vccd1 _3281_/X sky130_fd_sc_hd__mux2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _2227_/X _3539_/A _2232_/S vssd1 vssd1 vccd1 vccd1 _2234_/B sky130_fd_sc_hd__mux2_1
X_2163_ _1959_/C _2158_/X _2160_/X _2162_/X vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__a22o_1
X_2094_ _2094_/A _2189_/A vssd1 vssd1 vccd1 vccd1 _2094_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1948__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2996_ _3199_/B _2997_/C _2997_/A vssd1 vssd1 vccd1 vccd1 _2998_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1947_ _1947_/A vssd1 vssd1 vccd1 vccd1 _1948_/C sky130_fd_sc_hd__inv_2
X_1878_ _4083_/Q vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__inv_2
XFILLER_0_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2779__A _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3617_ _3635_/A0 hold183/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3617_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3548_ _3540_/A _3540_/B _3543_/B vssd1 vssd1 vccd1 vccd1 _3548_/X sky130_fd_sc_hd__o21ba_1
X_3479_ _3497_/A _3479_/B vssd1 vssd1 vccd1 vccd1 _4020_/D sky130_fd_sc_hd__and2_1
XANTENNA__2010__C _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2850_ _2674_/X _2835_/Y _2849_/X vssd1 vssd1 vccd1 vccd1 _3786_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2781_ _2813_/A _2781_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__and3_1
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold206 _3441_/X vssd1 vssd1 vccd1 vccd1 _3997_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold217 _3697_/Q vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _3635_/A0 hold191/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3402_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold228 _3380_/X vssd1 vssd1 vccd1 vccd1 _3948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _3945_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _2667_/X _3322_/X _3332_/X vssd1 vssd1 vccd1 vccd1 _3925_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _2661_/X _3257_/Y _3263_/X vssd1 vssd1 vccd1 vccd1 _3900_/D sky130_fd_sc_hd__a21o_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _2230_/A _2424_/B _2215_/C vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__or3_1
X_3195_ _3195_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3195_/X sky130_fd_sc_hd__or2_1
X_2146_ _2137_/X _2145_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3540_/B sky130_fd_sc_hd__mux2_2
X_2077_ _2075_/X _2076_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2077_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3395__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2979_ _3320_/A _2982_/B vssd1 vssd1 vccd1 vccd1 _2979_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold740 _4033_/Q vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout79_A _1863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3905_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2000_ _2153_/S _2614_/A _1998_/X _1987_/A vssd1 vssd1 vccd1 vccd1 _2194_/B sky130_fd_sc_hd__a22o_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3951_ _4105_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ _3834_/Q _3833_/Q _3830_/Q _3829_/Q vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__or4_2
X_3882_ _4092_/CLK _3882_/D vssd1 vssd1 vccd1 vccd1 _3882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2833_ _2834_/A _2834_/B vssd1 vssd1 vccd1 vccd1 _3358_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3377__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2764_ _2655_/X _2761_/X _2763_/X vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1945__B _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2695_ _2658_/X _2690_/Y _2694_/X vssd1 vssd1 vccd1 vccd1 _3722_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ hold669/X _2923_/B _3084_/Y _3123_/A vssd1 vssd1 vccd1 vccd1 _3316_/X sky130_fd_sc_hd__o211a_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3247_/A _3247_/B vssd1 vssd1 vccd1 vccd1 _3889_/D sky130_fd_sc_hd__or2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3301__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3178_ hold571/X _3189_/S _3177_/X _3497_/A vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__o211a_1
X_2129_ _2256_/A _2165_/B _3551_/A vssd1 vssd1 vccd1 vccd1 _2129_/X sky130_fd_sc_hd__and3_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold581 _4030_/Q vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 _3684_/X vssd1 vssd1 vccd1 vccd1 _3871_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _4100_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__buf_1
X_2480_ _3460_/A _2466_/X _2479_/X _2698_/A vssd1 vssd1 vccd1 vccd1 _3690_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2877__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3101_ _3099_/A _3060_/B _3036_/X _3100_/Y vssd1 vssd1 vccd1 vccd1 _3102_/D sky130_fd_sc_hd__a31oi_1
X_4081_ _4081_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
X_3032_ _3032_/A _3032_/B vssd1 vssd1 vccd1 vccd1 _3033_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ _3938_/CLK _3934_/D vssd1 vssd1 vccd1 vccd1 _3934_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2496__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3865_ _4072_/CLK _3865_/D vssd1 vssd1 vccd1 vccd1 _3865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2816_ _3640_/B _2854_/A vssd1 vssd1 vccd1 vccd1 _2831_/C sky130_fd_sc_hd__nand2_2
XANTENNA__1956__A _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3796_ _3803_/CLK _3796_/D vssd1 vssd1 vccd1 vccd1 _3796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2747_ _2658_/X _2742_/X _2746_/X vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2678_ _3566_/A _2382_/Y _2648_/Y _2677_/X vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__o31a_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2089__A0 _2119_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1866__A _3693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3860_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1980_ hold589/X _1890_/Y _1979_/X vssd1 vssd1 vccd1 vccd1 _2268_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3650_ _3654_/A _3650_/B _3656_/C vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3581_ _3581_/A _3596_/B vssd1 vssd1 vccd1 vccd1 _3581_/Y sky130_fd_sc_hd__nor2_1
X_2601_ _3637_/A0 hold179/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__mux2_1
X_2532_ _2355_/Y _2551_/B _2512_/A vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ _2232_/S _2461_/Y _3551_/B _2392_/A vssd1 vssd1 vccd1 vccd1 _2463_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3504__B1 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2394_ _2385_/A _2393_/X _2390_/Y vssd1 vssd1 vccd1 vccd1 _2394_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _4072_/CLK _4064_/D vssd1 vssd1 vccd1 vccd1 _4064_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2546__S _2588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3015_ _3857_/Q _3856_/Q _3032_/A vssd1 vssd1 vccd1 vccd1 _3027_/A sky130_fd_sc_hd__and3_1
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2469__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2794__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3917_ _4095_/CLK _3917_/D vssd1 vssd1 vccd1 vccd1 _3917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3848_ _4029_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_3779_ _3794_/CLK _3779_/D vssd1 vssd1 vccd1 vccd1 _3779_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout110 _3352_/A vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_8x305_116 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_116/HI io_out[24] sky130_fd_sc_hd__conb_1
XFILLER_0_75_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1963_ _3602_/A _2647_/A _1962_/X _1958_/X vssd1 vssd1 vccd1 vccd1 _1963_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2776__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3702_ _4072_/CLK _3702_/D vssd1 vssd1 vccd1 vccd1 _3702_/Q sky130_fd_sc_hd__dfxtp_1
X_1894_ _1895_/A _1895_/B vssd1 vssd1 vccd1 vccd1 _2616_/A sky130_fd_sc_hd__nand2_4
X_3633_ _3633_/A0 hold199/X _3639_/S vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3564_ _3564_/A _3564_/B vssd1 vssd1 vccd1 vccd1 _3564_/X sky130_fd_sc_hd__or2_1
X_3495_ _3497_/A _3495_/B vssd1 vssd1 vccd1 vccd1 _4028_/D sky130_fd_sc_hd__and2_1
X_2515_ _3973_/Q _4070_/Q _4062_/Q hold63/A _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2516_/B sky130_fd_sc_hd__mux4_1
X_2446_ _3946_/Q _3891_/Q _3697_/Q _4075_/Q _2584_/S0 _2584_/S1 vssd1 vssd1 vccd1
+ vccd1 _2447_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_75_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2377_ _2456_/B vssd1 vssd1 vccd1 vccd1 _2377_/Y sky130_fd_sc_hd__inv_2
X_4047_ _4047_/CLK _4047_/D vssd1 vssd1 vccd1 vccd1 _4047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2300_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2347_/S sky130_fd_sc_hd__inv_2
X_3280_ _3284_/A _3280_/B vssd1 vssd1 vccd1 vccd1 _3907_/D sky130_fd_sc_hd__and2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _3691_/Q _2230_/A _2226_/X _2230_/Y vssd1 vssd1 vccd1 vccd1 _3539_/A sky130_fd_sc_hd__a22o_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2885__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2162_ _2158_/S _2161_/X _2155_/S vssd1 vssd1 vccd1 vccd1 _2162_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2096__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2093_ _2238_/A _2093_/B vssd1 vssd1 vccd1 vccd1 _2189_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1948__B _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2749__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2995_ _2962_/A _2991_/X _2994_/Y vssd1 vssd1 vccd1 vccd1 _2995_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1946_ _2610_/A _1945_/Y _3602_/A vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__a21bo_1
X_1877_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3467_/A sky130_fd_sc_hd__inv_2
X_3616_ _1863_/Y hold235/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3616_/X sky130_fd_sc_hd__mux2_1
X_3547_ _1844_/A _3564_/B _3545_/Y _3546_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _4034_/D
+ sky130_fd_sc_hd__o221a_1
X_3478_ _1845_/A hold637/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3479_/B sky130_fd_sc_hd__mux2_1
X_2429_ _2571_/A _2571_/D vssd1 vssd1 vccd1 vccd1 _2430_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2795__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2780_ _3322_/A _2872_/A vssd1 vssd1 vccd1 vccd1 _2795_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2600__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 _4071_/Q vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _3965_/Q vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _3634_/A0 hold51/X _3406_/S vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__mux2_1
Xhold218 _2597_/X vssd1 vssd1 vccd1 vccd1 _3697_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3332_ _3654_/A _3332_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3332_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3269_/A _3263_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__and3_1
X_3194_ hold597/X _3189_/S _3193_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3194_/X sky130_fd_sc_hd__o211a_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2268_/A _2421_/A vssd1 vssd1 vccd1 vccd1 _2215_/C sky130_fd_sc_hd__nor2_1
X_2145_ _1959_/C _2140_/X _2142_/X _2144_/X vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2076_ _3931_/Q _3923_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2978_ _2984_/B _2978_/B vssd1 vssd1 vccd1 vccd1 _2982_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1929_ _1929_/A _1996_/S vssd1 vssd1 vccd1 vccd1 _1929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold730 _3694_/Q vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _4035_/Q vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2212__B _3551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__B1 _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ _4080_/CLK _3950_/D vssd1 vssd1 vccd1 vccd1 _3950_/Q sky130_fd_sc_hd__dfxtp_1
X_2901_ _3832_/Q _3831_/Q vssd1 vssd1 vccd1 vccd1 _3099_/C sky130_fd_sc_hd__or2_2
X_3881_ _4031_/CLK _3881_/D vssd1 vssd1 vccd1 vccd1 _3881_/Q sky130_fd_sc_hd__dfxtp_1
X_2832_ _2678_/X _2815_/X _2831_/X vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__a21o_1
X_2763_ _2813_/A _2763_/B _2777_/C vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2694_ _3269_/A _2694_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__and3_1
XFILLER_0_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3315_ _3320_/A _3315_/B vssd1 vssd1 vccd1 vccd1 _3919_/D sky130_fd_sc_hd__or2_1
X_3246_ _4042_/Q _1852_/A _3496_/S vssd1 vssd1 vccd1 vccd1 _3246_/X sky130_fd_sc_hd__mux2_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3177_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__or2_1
X_2128_ _2119_/X _2127_/X _2164_/S vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__mux2_2
X_2059_ _2057_/X _2058_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2059_/X sky130_fd_sc_hd__mux2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2576__C1 _2612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 _4019_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__buf_1
XANTENNA_fanout91_A _3467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 _2683_/X vssd1 vssd1 vccd1 vccd1 _3717_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _3473_/X vssd1 vssd1 vccd1 vccd1 _4017_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _3669_/X vssd1 vssd1 vccd1 vccd1 _4100_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3100_ _3100_/A _3285_/B _3100_/C vssd1 vssd1 vccd1 vccd1 _3100_/Y sky130_fd_sc_hd__nor3_1
X_4080_ _4080_/CLK hold90/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
X_3031_ _3854_/Q _3054_/A _3855_/Q vssd1 vssd1 vccd1 vccd1 _3032_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3295__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3933_ _4088_/CLK _3933_/D vssd1 vssd1 vccd1 vccd1 _3933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4072_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2270__B2 _1867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3864_ _4072_/CLK _3864_/D vssd1 vssd1 vccd1 vccd1 _3864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ _3640_/B _2854_/A vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__and2_2
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3795_ _3795_/CLK _3795_/D vssd1 vssd1 vccd1 vccd1 _3795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2746_ _2805_/A _2746_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2746_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2677_ _2677_/A _2677_/B vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3497_/A _3229_/B vssd1 vssd1 vccd1 vccd1 _3880_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3286__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold390 _3773_/Q vssd1 vssd1 vccd1 vccd1 _2819_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3277__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3580_ _2642_/A _2646_/D _3579_/X _3227_/A vssd1 vssd1 vccd1 vccd1 _3580_/X sky130_fd_sc_hd__o211a_1
X_2600_ _3636_/A0 hold241/X _2603_/S vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__mux2_1
X_2531_ _2573_/S _3518_/A _2529_/X _2530_/Y vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__o22a_1
X_2462_ _2573_/S _2461_/Y _3551_/B vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2099__S _2159_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3504__A1 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2393_ _2512_/A _2393_/B _2551_/B vssd1 vssd1 vccd1 vccd1 _2393_/X sky130_fd_sc_hd__or3_2
X_4063_ _4081_/CLK _4063_/D vssd1 vssd1 vccd1 vccd1 _4063_/Q sky130_fd_sc_hd__dfxtp_1
X_3014_ _3855_/Q _3854_/Q _3054_/A vssd1 vssd1 vccd1 vccd1 _3032_/A sky130_fd_sc_hd__and3_1
XANTENNA__3440__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3916_ _4095_/CLK _3916_/D vssd1 vssd1 vccd1 vccd1 _3916_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2243__A1 _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3847_ _3862_/CLK _3847_/D vssd1 vssd1 vccd1 vccd1 _3847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _3778_/CLK _3778_/D vssd1 vssd1 vccd1 vccd1 _3778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2729_ _2421_/A _2728_/X _2734_/S vssd1 vssd1 vccd1 vccd1 _2729_/X sky130_fd_sc_hd__mux2_1
Xfanout111 _3352_/A vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__clkbuf_4
Xfanout100 _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3687_/C1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3431__A0 _3635_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1993__A0 _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwrapped_8x305_117 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_117/HI io_out[25] sky130_fd_sc_hd__conb_1
XANTENNA_output35_A _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3422__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1962_ _3321_/A _3321_/B _3340_/A _2296_/B vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3701_ _4080_/CLK _3701_/D vssd1 vssd1 vccd1 vccd1 _3701_/Q sky130_fd_sc_hd__dfxtp_1
X_1893_ _2008_/C _3600_/B _3907_/Q vssd1 vssd1 vccd1 vccd1 _1895_/B sky130_fd_sc_hd__or3_4
XFILLER_0_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3632_ _3676_/A0 hold175/X _3639_/S vssd1 vssd1 vccd1 vccd1 _3632_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3563_ _3554_/Y _3561_/Y _3562_/X _3554_/B hold679/X vssd1 vssd1 vccd1 vccd1 _3563_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3507__A _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2514_ _2392_/X _2508_/C _2391_/X vssd1 vssd1 vccd1 vccd1 _2514_/Y sky130_fd_sc_hd__a21oi_1
X_3494_ hold694/X _4028_/Q _3494_/S vssd1 vssd1 vccd1 vccd1 _3494_/X sky130_fd_sc_hd__mux2_1
X_2445_ _2585_/A _2445_/B vssd1 vssd1 vccd1 vccd1 _2445_/Y sky130_fd_sc_hd__nand2b_1
X_2376_ _2376_/A _2376_/B _2376_/C vssd1 vssd1 vccd1 vccd1 _2456_/B sky130_fd_sc_hd__and3_1
X_4046_ _4047_/CLK _4046_/D vssd1 vssd1 vccd1 vccd1 _4046_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3661__A0 _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3413__A0 _3636_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2216__A1 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3404__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2230_/A _2230_/B vssd1 vssd1 vccd1 vccd1 _2230_/Y sky130_fd_sc_hd__nor2_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3062__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2161_ _3904_/Q _3786_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2161_/X sky130_fd_sc_hd__mux2_1
X_2092_ _2220_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2094_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2994_ _2962_/A _2991_/X _3114_/A vssd1 vssd1 vccd1 vccd1 _2994_/Y sky130_fd_sc_hd__o21ai_1
X_1945_ _2616_/A _2180_/B vssd1 vssd1 vccd1 vccd1 _1945_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_9_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1876_ _2891_/A vssd1 vssd1 vccd1 vccd1 _2986_/A sky130_fd_sc_hd__inv_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3615_ _3633_/A0 hold245/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3615_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3546_ _2621_/A _3554_/B hold368/X vssd1 vssd1 vccd1 vccd1 _3546_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout104_A _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3477_ _3497_/A _3477_/B vssd1 vssd1 vccd1 vccd1 _4019_/D sky130_fd_sc_hd__and2_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2428_ _2362_/S _2355_/Y _2349_/X _2347_/S vssd1 vssd1 vccd1 vccd1 _2428_/X sky130_fd_sc_hd__a211o_1
X_2359_ _2260_/X _2283_/X _2356_/Y _2181_/Y vssd1 vssd1 vccd1 vccd1 _2360_/B sky130_fd_sc_hd__a31o_1
X_4029_ _4029_/CLK _4029_/D vssd1 vssd1 vccd1 vccd1 _4029_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3634__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3625__A0 _1863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold208 _3628_/X vssd1 vssd1 vccd1 vccd1 _4071_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _3633_/A0 hold147/X _3406_/S vssd1 vssd1 vccd1 vccd1 _3400_/X sky130_fd_sc_hd__mux2_1
Xhold219 _4066_/Q vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_3331_ _2664_/X _3322_/X _3330_/X vssd1 vssd1 vccd1 vccd1 _3924_/D sky130_fd_sc_hd__a21o_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _2658_/X _3257_/Y _3261_/X vssd1 vssd1 vccd1 vccd1 _3899_/D sky130_fd_sc_hd__a21o_1
X_3193_ _3193_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__or2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2256_/A _2211_/Y _2212_/Y _2573_/S vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__a211o_1
X_2144_ _2158_/S _2143_/X _2155_/S vssd1 vssd1 vccd1 vccd1 _2144_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_15_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3616__A0 _1863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2075_ _4084_/Q _3939_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1959__B _2158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2977_ _2978_/B _3131_/A _2977_/C vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1928_ _1988_/A _2180_/B _3596_/A vssd1 vssd1 vccd1 vccd1 _2227_/S sky130_fd_sc_hd__a21oi_4
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ _3880_/Q vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__inv_2
Xhold720 _4028_/Q vssd1 vssd1 vccd1 vccd1 _3048_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _3694_/Q vssd1 vssd1 vccd1 vccd1 _3468_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _4036_/Q vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _3529_/A _3529_/B vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3607__A0 _3634_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4045_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2830__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2346__A0 _3507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__A1 _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2655__S _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2900_ _3199_/B _2988_/B vssd1 vssd1 vccd1 vccd1 _3275_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3880_ _4092_/CLK _3880_/D vssd1 vssd1 vccd1 vccd1 _3880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2831_ _2869_/A _2831_/B _2831_/C vssd1 vssd1 vccd1 vccd1 _2831_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2762_ _3322_/A _2854_/A vssd1 vssd1 vccd1 vccd1 _2777_/C sky130_fd_sc_hd__nand2_2
X_2693_ _2655_/X _2690_/Y _2692_/X vssd1 vssd1 vccd1 vccd1 _2693_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2888__A1 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ hold707/X _3313_/X _3314_/S vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__mux2_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3247_/A _3245_/B vssd1 vssd1 vccd1 vccd1 _3888_/D sky130_fd_sc_hd__or2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3247_/A _3176_/B vssd1 vssd1 vccd1 vccd1 _3850_/D sky130_fd_sc_hd__or2_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2127_ _1959_/C _2122_/X _2124_/X _2126_/X vssd1 vssd1 vccd1 vccd1 _2127_/X sky130_fd_sc_hd__a22o_1
X_2058_ _3932_/Q _3924_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__mux2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2812__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold561 _3858_/Q vssd1 vssd1 vccd1 vccd1 _3191_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _3189_/X vssd1 vssd1 vccd1 vccd1 _3190_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _3820_/Q vssd1 vssd1 vccd1 vccd1 _2982_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _3811_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _3798_/Q vssd1 vssd1 vccd1 vccd1 _2877_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3030_ _4024_/Q _3030_/B vssd1 vssd1 vccd1 vccd1 _3055_/A sky130_fd_sc_hd__xnor2_1
X_3932_ _3938_/CLK _3932_/D vssd1 vssd1 vccd1 vccd1 _3932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ _4072_/CLK _3863_/D vssd1 vssd1 vccd1 vccd1 _3863_/Q sky130_fd_sc_hd__dfxtp_1
X_2814_ _2678_/X _2797_/X _2813_/X vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3794_ _3794_/CLK _3794_/D vssd1 vssd1 vccd1 vccd1 _3794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2745_ _2655_/X _2742_/X _2744_/X vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__a21o_1
X_2676_ _2813_/A _2676_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _1846_/Y _1859_/Y _3494_/S vssd1 vssd1 vccd1 vccd1 _3228_/X sky130_fd_sc_hd__mux2_1
X_3159_ _3165_/B _3159_/B vssd1 vssd1 vccd1 vccd1 _3159_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3210__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 _3165_/X vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _2820_/X vssd1 vssd1 vccd1 vccd1 _3773_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2530_ _3637_/A0 _2529_/B _2573_/S vssd1 vssd1 vccd1 vccd1 _2530_/Y sky130_fd_sc_hd__o21ai_1
X_2461_ _3634_/A0 _2458_/X _2460_/X vssd1 vssd1 vccd1 vccd1 _2461_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2392_ _2392_/A _2612_/B _2511_/S vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__and3_1
X_4062_ _4073_/CLK _4062_/D vssd1 vssd1 vccd1 vccd1 _4062_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3268__A1 _2667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3013_ _3853_/Q _3852_/Q _3043_/A vssd1 vssd1 vccd1 vccd1 _3054_/A sky130_fd_sc_hd__and3_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3915_ _4092_/CLK _3915_/D vssd1 vssd1 vccd1 vccd1 _3915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3846_ _3846_/CLK _3846_/D vssd1 vssd1 vccd1 vccd1 _3846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3777_ _3794_/CLK _3777_/D vssd1 vssd1 vccd1 vccd1 _3777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2728_ _3558_/B _2733_/S _2727_/X vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__2951__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2659_ _2652_/Y _2658_/X _2657_/X vssd1 vssd1 vccd1 vccd1 _3710_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout112 _2698_/A vssd1 vssd1 vccd1 vccd1 _3352_/A sky130_fd_sc_hd__clkbuf_2
Xfanout101 _2953_/B1 vssd1 vssd1 vccd1 vccd1 _3471_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwrapped_8x305_118 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_118/HI io_out[26] sky130_fd_sc_hd__conb_1
X_3700_ _4081_/CLK _3700_/D vssd1 vssd1 vccd1 vccd1 _3700_/Q sky130_fd_sc_hd__dfxtp_1
X_1961_ _2834_/A _2834_/B vssd1 vssd1 vccd1 vccd1 _3341_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1892_ _2008_/C _3600_/B _2737_/A vssd1 vssd1 vccd1 vccd1 _1895_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3631_ _3631_/A _3631_/B vssd1 vssd1 vccd1 vccd1 _3639_/S sky130_fd_sc_hd__or2_4
X_3562_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3562_/X sky130_fd_sc_hd__or2_1
X_2513_ _2392_/A _2510_/X _2512_/X _2612_/B vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__o211a_1
X_3493_ _3497_/A _3493_/B vssd1 vssd1 vccd1 vccd1 _4027_/D sky130_fd_sc_hd__and2_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2444_ _3978_/Q hold59/A _3962_/Q _3954_/Q _2582_/S0 _2582_/S1 vssd1 vssd1 vccd1
+ vccd1 _2445_/B sky130_fd_sc_hd__mux4_1
X_2375_ _2424_/B _2374_/Y _2484_/A _2372_/Y vssd1 vssd1 vccd1 vccd1 _2375_/X sky130_fd_sc_hd__a2bb2o_1
X_4045_ _4045_/CLK _4045_/D vssd1 vssd1 vccd1 vccd1 _4045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3829_ _4095_/CLK _3829_/D vssd1 vssd1 vccd1 vccd1 _3829_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1975__A1 _3322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2658__S _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _2160_/A _2160_/B vssd1 vssd1 vccd1 vccd1 _2160_/X sky130_fd_sc_hd__or2_1
X_2091_ _1988_/A _2089_/X _2614_/A _2119_/S vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__a2bb2o_2
XANTENNA__3643__A1 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2993_ _2991_/X hold648/X _3114_/A vssd1 vssd1 vccd1 vccd1 _2993_/Y sky130_fd_sc_hd__o21ai_1
X_1944_ _3602_/A _3201_/A vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__and2_1
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1875_ _2992_/A vssd1 vssd1 vccd1 vccd1 _2969_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3518__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _3676_/A0 hold263/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3614_/X sky130_fd_sc_hd__mux2_1
X_3545_ _3554_/B _3545_/B vssd1 vssd1 vccd1 vccd1 _3545_/Y sky130_fd_sc_hd__nor2_1
X_3476_ _1846_/A hold571/X _3494_/S vssd1 vssd1 vccd1 vccd1 _3477_/B sky130_fd_sc_hd__mux2_1
X_2427_ _2571_/A _2427_/B vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__or2_1
X_2358_ _2260_/X _2283_/X _2356_/Y vssd1 vssd1 vccd1 vccd1 _2360_/A sky130_fd_sc_hd__a21oi_1
X_2289_ _2289_/A vssd1 vssd1 vccd1 vccd1 _2289_/Y sky130_fd_sc_hd__inv_2
X_4028_ _4092_/CLK _4028_/D vssd1 vssd1 vccd1 vccd1 _4028_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3399__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3389__A0 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold209 _4069_/Q vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
X_3330_ _3654_/A _3330_/B _3338_/C vssd1 vssd1 vccd1 vccd1 _3330_/X sky130_fd_sc_hd__and3_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3269_/A _3261_/B _3273_/C vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__and3_1
X_3192_ hold729/X _3189_/S _3191_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__o211a_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2256_/A _3551_/A vssd1 vssd1 vccd1 vccd1 _2212_/Y sky130_fd_sc_hd__nor2_1
X_2143_ _3902_/Q _3784_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__mux2_1
X_2074_ _2070_/X _2073_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2074_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1959__C _1959_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2976_ _3199_/A _2976_/B _3817_/Q vssd1 vssd1 vccd1 vccd1 _2978_/B sky130_fd_sc_hd__and3_1
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1927_ hold636/X _1890_/Y _1925_/X vssd1 vssd1 vccd1 vccd1 _3540_/A sky130_fd_sc_hd__o21a_4
X_1858_ _3881_/Q vssd1 vssd1 vccd1 vccd1 _1858_/Y sky130_fd_sc_hd__inv_2
Xhold710 _3065_/Y vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _3057_/X vssd1 vssd1 vccd1 vccd1 _3058_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3682__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold743 _4034_/Q vssd1 vssd1 vccd1 vccd1 hold743/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 _3706_/Q vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
X_3528_ _3528_/A _3528_/B vssd1 vssd1 vccd1 vccd1 _3528_/Y sky130_fd_sc_hd__xnor2_1
X_3459_ hold728/X _3470_/B hold280/X _3471_/C1 vssd1 vssd1 vccd1 vccd1 _3459_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2327__A _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ _2674_/X _2815_/X _2829_/X vssd1 vssd1 vccd1 vccd1 _3778_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2761_ _3322_/A _2854_/A vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__and2_2
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2692_ _2869_/A _2692_/B _2706_/C vssd1 vssd1 vccd1 vccd1 _2692_/X sky130_fd_sc_hd__and3_1
XANTENNA_1 _3683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _2988_/B _3312_/X _3120_/Y vssd1 vssd1 vccd1 vccd1 _3313_/X sky130_fd_sc_hd__a21o_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _4041_/Q _1853_/A _3494_/S vssd1 vssd1 vccd1 vccd1 _3244_/X sky130_fd_sc_hd__mux2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _4018_/Q hold681/X _3189_/S vssd1 vssd1 vccd1 vccd1 _3175_/X sky130_fd_sc_hd__mux2_1
X_2126_ _2151_/S _2125_/X _2155_/S vssd1 vssd1 vccd1 vccd1 _2126_/X sky130_fd_sc_hd__o21a_1
X_2057_ _4085_/Q _3940_/Q _2157_/S vssd1 vssd1 vccd1 vccd1 _2057_/X sky130_fd_sc_hd__mux2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3677__S _3683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2959_ _2962_/A _2992_/A vssd1 vssd1 vccd1 vccd1 _2997_/C sky130_fd_sc_hd__and2_1
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold551 hold737/X vssd1 vssd1 vccd1 vccd1 _1841_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold562 _3192_/X vssd1 vssd1 vccd1 vccd1 _3858_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _3825_/Q vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold584 _2946_/Y vssd1 vssd1 vccd1 vccd1 _3811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _2986_/B vssd1 vssd1 vccd1 vccd1 _2983_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _3860_/Q vssd1 vssd1 vccd1 vccd1 _3195_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3461__C1 _3471_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3931_ _3939_/CLK _3931_/D vssd1 vssd1 vccd1 vccd1 _3931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3862_ _3862_/CLK _3862_/D vssd1 vssd1 vccd1 vccd1 _3862_/Q sky130_fd_sc_hd__dfxtp_1
X_2813_ _2813_/A _2813_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3793_ _3794_/CLK _3793_/D vssd1 vssd1 vccd1 vccd1 _3793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2744_ _2813_/A _2744_/B _2758_/C vssd1 vssd1 vccd1 vccd1 _2744_/X sky130_fd_sc_hd__and3_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2675_ _2652_/Y _2674_/X _2673_/X vssd1 vssd1 vccd1 vccd1 _3715_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _3227_/A _3227_/B vssd1 vssd1 vccd1 vccd1 _3879_/D sky130_fd_sc_hd__nand2_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ hold292/X _3199_/B _3157_/X vssd1 vssd1 vccd1 vccd1 _3159_/B sky130_fd_sc_hd__o21ai_1
X_2109_ _1959_/C _2104_/X _2106_/X _2108_/X vssd1 vssd1 vccd1 vccd1 _2109_/X sky130_fd_sc_hd__a22o_1
X_3089_ _2988_/B _3057_/X _3081_/Y _3136_/A _3087_/Y vssd1 vssd1 vccd1 vccd1 _3089_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold381 _3166_/X vssd1 vssd1 vccd1 vccd1 _3846_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _3778_/Q vssd1 vssd1 vccd1 vccd1 _2829_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2721__A1 _3551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 _3756_/Q vssd1 vssd1 vccd1 vccd1 _2781_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2580__S0 _2584_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2788__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2460_ _2508_/A _2453_/Y _2454_/Y _2458_/X _2459_/X vssd1 vssd1 vccd1 vccd1 _2460_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2399__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2391_ _2009_/A _1977_/B _2008_/C _2009_/B vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _4081_/CLK _4061_/D vssd1 vssd1 vccd1 vccd1 _4061_/Q sky130_fd_sc_hd__dfxtp_1
X_3012_ _3852_/Q _3043_/A vssd1 vssd1 vccd1 vccd1 _3040_/A sky130_fd_sc_hd__and2_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3914_ _4095_/CLK _3914_/D vssd1 vssd1 vccd1 vccd1 _3914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3845_ _3846_/CLK _3845_/D vssd1 vssd1 vccd1 vccd1 _3845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ _3791_/CLK _3776_/D vssd1 vssd1 vccd1 vccd1 _3776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2727_ _2733_/S _2732_/B _2727_/C vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__or3_1
XFILLER_0_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2160__A _2160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2658_ _2551_/A _2553_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__mux2_8
X_2589_ _2393_/B _2588_/X _2577_/X vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout113 input23/X vssd1 vssd1 vccd1 vccd1 _2698_/A sky130_fd_sc_hd__buf_4
XANTENNA__2703__A1 _2671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 input23/X vssd1 vssd1 vccd1 vccd1 _2953_/B1 sky130_fd_sc_hd__buf_2
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2942__A1 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_8x305_119 vssd1 vssd1 vccd1 vccd1 wrapped_8x305_119/HI io_out[27] sky130_fd_sc_hd__conb_1
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ _2834_/A _2834_/B vssd1 vssd1 vccd1 vccd1 _3340_/A sky130_fd_sc_hd__and2_2
X_1891_ _3602_/A _3600_/B vssd1 vssd1 vccd1 vccd1 _1996_/S sky130_fd_sc_hd__or2_4
X_3630_ _3639_/A0 hold261/X _3630_/S vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__mux2_1
X_3561_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3561_/Y sky130_fd_sc_hd__nand2_1
X_2512_ _2512_/A _2512_/B vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3492_ _3575_/A hold597/X _3494_/S vssd1 vssd1 vccd1 vccd1 _3493_/B sky130_fd_sc_hd__mux2_1
X_2443_ _2585_/A _2442_/X _3720_/Q vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__a21oi_1
X_2374_ _2268_/A _2378_/C _2484_/A vssd1 vssd1 vccd1 vccd1 _2374_/Y sky130_fd_sc_hd__o21bai_1
X_4113_ _4113_/CLK _4113_/D vssd1 vssd1 vccd1 vccd1 _4113_/Q sky130_fd_sc_hd__dfxtp_1
X_4044_ _4101_/CLK _4044_/D vssd1 vssd1 vccd1 vccd1 _4044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3828_ _4077_/CLK _3828_/D vssd1 vssd1 vccd1 vccd1 _3828_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1975__A2 _2296_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3759_ _3767_/CLK _3759_/D vssd1 vssd1 vccd1 vccd1 _3759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output40_A _3808_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ _1959_/C _1988_/Y _2089_/X _1988_/A vssd1 vssd1 vccd1 vccd1 _2093_/B sky130_fd_sc_hd__o22a_4
XANTENNA__2674__S _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2992_ _2992_/A _3004_/A vssd1 vssd1 vccd1 vccd1 _2992_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2603__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1943_ _3322_/A _2296_/B _3321_/A _1943_/D vssd1 vssd1 vccd1 vccd1 _3201_/A sky130_fd_sc_hd__and4_4
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1874_ _2960_/A vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__inv_2
X_3613_ _3874_/Q _3873_/Q _3613_/C vssd1 vssd1 vccd1 vccd1 _3621_/S sky130_fd_sc_hd__or3_4
XFILLER_0_71_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3544_ _3539_/Y _3543_/Y _3544_/S vssd1 vssd1 vccd1 vccd1 _3545_/B sky130_fd_sc_hd__mux2_1
X_3475_ _3587_/A _3475_/B vssd1 vssd1 vccd1 vccd1 _4018_/D sky130_fd_sc_hd__and2_1
X_2426_ _2423_/X _2528_/B _2570_/A vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3331__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2357_ _1945_/Y _2247_/X _2356_/Y _2616_/A _2181_/Y vssd1 vssd1 vccd1 vccd1 _2357_/X
+ sky130_fd_sc_hd__o221a_1
X_2288_ _2288_/A _2288_/B vssd1 vssd1 vccd1 vccd1 _2289_/A sky130_fd_sc_hd__nor2_1
XANTENNA__2517__S0 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4027_ _4092_/CLK _4027_/D vssd1 vssd1 vccd1 vccd1 _4027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _2655_/X _3257_/Y _3259_/X vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__a21o_1
X_3191_ _3191_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3191_/X sky130_fd_sc_hd__or2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2189_/A _2209_/X _2210_/X vssd1 vssd1 vccd1 vccd1 _2211_/Y sky130_fd_sc_hd__a21oi_1
X_2142_ _2142_/A _2142_/B vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__or2_1
X_2073_ _2071_/X _2072_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__mux2_1
X_2975_ _3199_/A _3817_/Q _2974_/X _2976_/B vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3529__A _3529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1926_ _4094_/Q _1890_/Y _1925_/X vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1857_ _3882_/Q vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__inv_2
Xhold700 _2890_/Y vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 _3068_/X vssd1 vssd1 vccd1 vccd1 _3832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _4029_/Q vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 _3705_/Q vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 _3059_/X vssd1 vssd1 vccd1 vccd1 _3829_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ _3518_/A _3518_/B _3526_/X vssd1 vssd1 vccd1 vccd1 _3528_/B sky130_fd_sc_hd__a21oi_1
X_3458_ _3458_/A _3470_/B vssd1 vssd1 vccd1 vccd1 _3458_/Y sky130_fd_sc_hd__nand2_1
X_2409_ _2409_/A _2409_/B vssd1 vssd1 vccd1 vccd1 _2940_/B sky130_fd_sc_hd__nor2_1
X_3389_ _3676_/A0 hold75/X _3396_/S vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2351__A1_N _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4077_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2760_ _3321_/A _3321_/B _3640_/A vssd1 vssd1 vccd1 vccd1 _2854_/A sky130_fd_sc_hd__and3_2
X_2691_ _3323_/A _3258_/A vssd1 vssd1 vccd1 vccd1 _2706_/C sky130_fd_sc_hd__or2_2
XANTENNA_2 _3960_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ hold645/X _3125_/Y _3311_/X _3097_/Y vssd1 vssd1 vccd1 vccd1 _3312_/X sky130_fd_sc_hd__a211o_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3587_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3887_/D sky130_fd_sc_hd__nand2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3247_/A _3174_/B vssd1 vssd1 vccd1 vccd1 _3849_/D sky130_fd_sc_hd__or2_1
X_2125_ _3903_/Q _3785_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2052_/X _2055_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2056_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2958_ _2960_/A _3824_/Q vssd1 vssd1 vccd1 vccd1 _3120_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ _4099_/Q _1890_/Y _1907_/X vssd1 vssd1 vccd1 vccd1 _2160_/A sky130_fd_sc_hd__o21ai_4
X_2889_ _2982_/A _2984_/B vssd1 vssd1 vccd1 vccd1 _2974_/B sky130_fd_sc_hd__or2_1
Xhold530 _3752_/Q vssd1 vssd1 vccd1 vccd1 _2771_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _3238_/X vssd1 vssd1 vccd1 vccd1 _3239_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _2999_/Y vssd1 vssd1 vccd1 vccd1 _3825_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _4101_/Q vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2610__B _2737_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 _2983_/X vssd1 vssd1 vccd1 vccd1 _3820_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _3196_/X vssd1 vssd1 vccd1 vccd1 _3860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _3780_/Q vssd1 vssd1 vccd1 vccd1 _2837_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold536_A _3812_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3516__A1 _3506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput50 _3676_/A0 vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XANTENNA__3452__A0 _1867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _3939_/CLK _3930_/D vssd1 vssd1 vccd1 vccd1 _3930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3861_ _4029_/CLK _3861_/D vssd1 vssd1 vccd1 vccd1 _3861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3792_ _3794_/CLK _3792_/D vssd1 vssd1 vccd1 vccd1 _3792_/Q sky130_fd_sc_hd__dfxtp_1
X_2812_ _2674_/X _2797_/X _2811_/X vssd1 vssd1 vccd1 vccd1 _3770_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2743_ _3340_/A _2872_/A vssd1 vssd1 vccd1 vccd1 _2758_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2674_ _2435_/A _2434_/X _2677_/B vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__mux2_8
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _1847_/Y _1860_/Y _3496_/S vssd1 vssd1 vccd1 vccd1 _3226_/X sky130_fd_sc_hd__mux2_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3157_ _3157_/A _3157_/B vssd1 vssd1 vccd1 vccd1 _3157_/X sky130_fd_sc_hd__or2_1
X_2108_ _2158_/S _2107_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2108_/X sky130_fd_sc_hd__o21a_1
X_3088_ _3088_/A _3088_/B vssd1 vssd1 vccd1 vccd1 _3090_/B sky130_fd_sc_hd__or2_1
XFILLER_0_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3443__A0 _1867_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2039_ _4082_/Q _3937_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2039_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold371 _3714_/Q vssd1 vssd1 vccd1 vccd1 _2669_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _3867_/Q vssd1 vssd1 vccd1 vccd1 _2408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _2782_/X vssd1 vssd1 vccd1 vccd1 _3756_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _3936_/Q vssd1 vssd1 vccd1 vccd1 _3356_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3682__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2580__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3434__A0 _3682_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2399__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2390_ _2009_/A _1977_/B _3602_/A _2009_/B vssd1 vssd1 vccd1 vccd1 _2390_/Y sky130_fd_sc_hd__a211oi_2
XANTENNA__2173__B1 _3676_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ _4073_/CLK _4060_/D vssd1 vssd1 vccd1 vccd1 _4060_/Q sky130_fd_sc_hd__dfxtp_1
X_3011_ _3851_/Q _3850_/Q _3849_/Q vssd1 vssd1 vccd1 vccd1 _3043_/A sky130_fd_sc_hd__and3_1
XANTENNA__3673__A0 _2180_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3425__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2706__A _2813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3913_ _4101_/CLK _3913_/D vssd1 vssd1 vccd1 vccd1 _3913_/Q sky130_fd_sc_hd__dfxtp_1
X_3844_ _3846_/CLK _3844_/D vssd1 vssd1 vccd1 vccd1 _3844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3775_ _3791_/CLK _3775_/D vssd1 vssd1 vccd1 vccd1 _3775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2726_ _3737_/Q _2726_/B vssd1 vssd1 vccd1 vccd1 _2727_/C sky130_fd_sc_hd__nor2_1
XANTENNA__2951__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2657_ _3269_/A _2657_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2588_ _2587_/X input8/X _2588_/S vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__mux2_1
Xfanout103 _2887_/A vssd1 vssd1 vccd1 vccd1 _3227_/A sky130_fd_sc_hd__buf_4
X_3209_ _3692_/Q _3201_/Y _3208_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3209_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3416__A0 _3639_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2616__A _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2942__A2 _2940_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 _2598_/X vssd1 vssd1 vccd1 vccd1 _3698_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1969__B1 _3540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1890_ _3602_/A _3600_/B vssd1 vssd1 vccd1 vccd1 _1890_/Y sky130_fd_sc_hd__nor2_8
X_3560_ _3553_/A _3550_/Y _3552_/B vssd1 vssd1 vccd1 vccd1 _3562_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2511_ _2361_/X _2508_/Y _2511_/S vssd1 vssd1 vccd1 vccd1 _2512_/B sky130_fd_sc_hd__mux2_1
X_3491_ _3497_/A _3491_/B vssd1 vssd1 vccd1 vccd1 _4026_/D sky130_fd_sc_hd__and2_1
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2442_ hold33/A _3994_/Q _4010_/Q _3986_/Q _2582_/S1 _2582_/S0 vssd1 vssd1 vccd1
+ vccd1 _2442_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2697__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2373_ _2424_/A _2373_/B vssd1 vssd1 vccd1 vccd1 _2378_/C sky130_fd_sc_hd__nor2_1
X_4112_ _4112_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
X_4043_ _4101_/CLK _4043_/D vssd1 vssd1 vccd1 vccd1 _4043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3827_ _4077_/CLK _3827_/D vssd1 vssd1 vccd1 vccd1 _3827_/Q sky130_fd_sc_hd__dfxtp_1
X_3758_ _3767_/CLK _3758_/D vssd1 vssd1 vccd1 vccd1 _3758_/Q sky130_fd_sc_hd__dfxtp_1
X_2709_ _2834_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _3640_/B sky130_fd_sc_hd__nor2_2
X_3689_ _3690_/CLK _3689_/D vssd1 vssd1 vccd1 vccd1 _3689_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3637__A0 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2860__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2471__S0 _2584_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2020__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2991_ _2992_/A _2990_/X _3004_/A vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _2230_/A _1942_/B vssd1 vssd1 vccd1 vccd1 _1943_/D sky130_fd_sc_hd__or2_1
X_1873_ _2990_/D vssd1 vssd1 vccd1 vccd1 _3106_/A sky130_fd_sc_hd__inv_2
XFILLER_0_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3612_ _3639_/A0 hold193/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3612_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_leaf_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3543_ _3543_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3543_/Y sky130_fd_sc_hd__xnor2_1
X_3474_ hold665/X hold723/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3475_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ _2424_/X _2484_/B _2484_/A vssd1 vssd1 vccd1 vccd1 _2528_/B sky130_fd_sc_hd__mux2_1
X_2356_ _4085_/Q _2356_/B vssd1 vssd1 vccd1 vccd1 _2356_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2287_ _2235_/Y _2246_/Y _2284_/X _2288_/B _2233_/X vssd1 vssd1 vccd1 vccd1 _2287_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3550__A _3551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2517__S1 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4026_ _4029_/CLK _4026_/D vssd1 vssd1 vccd1 vccd1 _4026_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2842__A1 _2661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2105__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3460__A _3460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2597__A0 _3633_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2015__S _2151_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2444__S0 _2582_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2222_/A _2049_/X _2094_/Y _2207_/X _2093_/B vssd1 vssd1 vccd1 vccd1 _2210_/X
+ sky130_fd_sc_hd__a32o_1
X_3190_ _3320_/A _3190_/B vssd1 vssd1 vccd1 vccd1 _3857_/D sky130_fd_sc_hd__or2_1
XFILLER_0_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2141_ _3713_/Q _3725_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2142_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2072_ _3774_/Q _3790_/Q _2152_/S vssd1 vssd1 vccd1 vccd1 _2072_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2824__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2974_ _2986_/A _2974_/B vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _4111_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1925_ _3602_/A _3600_/B _1925_/C vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__or3_2
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1856_ _3883_/Q vssd1 vssd1 vccd1 vccd1 _1856_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold712 _3837_/Q vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold701 _3833_/Q vssd1 vssd1 vccd1 vccd1 _2935_/B sky130_fd_sc_hd__buf_1
Xhold723 _4018_/Q vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 _3704_/Q vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _4032_/Q vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
X_3526_ _3518_/A _3518_/B _3520_/B vssd1 vssd1 vccd1 vccd1 _3526_/X sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout102_A input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3457_ _3467_/A _3457_/B vssd1 vssd1 vccd1 vccd1 _4009_/D sky130_fd_sc_hd__or2_1
X_2408_ _2408_/A _2408_/B _2408_/C _2408_/D vssd1 vssd1 vccd1 vccd1 _2409_/B sky130_fd_sc_hd__or4_1
X_3388_ _3604_/C _3675_/A vssd1 vssd1 vccd1 vccd1 _3396_/S sky130_fd_sc_hd__or2_4
X_2339_ _2345_/S _2338_/B _2181_/Y vssd1 vssd1 vccd1 vccd1 _2339_/Y sky130_fd_sc_hd__a21oi_1
X_4009_ _4014_/CLK _4009_/D vssd1 vssd1 vccd1 vccd1 _4009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3190__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2806__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2690_ _3323_/A _3258_/A vssd1 vssd1 vccd1 vccd1 _2690_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 hold499/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3311_ _3024_/A _3124_/Y _3304_/Y _4018_/Q vssd1 vssd1 vccd1 vccd1 _3311_/X sky130_fd_sc_hd__a22o_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _1839_/Y _1854_/Y _3494_/S vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__mux2_1
X_3173_ hold659/X _3849_/Q _3189_/S vssd1 vssd1 vccd1 vccd1 _3173_/X sky130_fd_sc_hd__mux2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2142_/A _2124_/B vssd1 vssd1 vccd1 vccd1 _2124_/X sky130_fd_sc_hd__or2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2053_/X _2054_/X _2142_/A vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2957_ _3199_/A _3199_/B vssd1 vssd1 vccd1 vccd1 _2957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1908_ _3911_/Q hold565/X _1996_/S vssd1 vssd1 vccd1 vccd1 _1908_/X sky130_fd_sc_hd__mux2_1
X_2888_ _2678_/X _2871_/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__a21o_1
X_1839_ _3575_/A vssd1 vssd1 vccd1 vccd1 _1839_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold520 _3694_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__clkbuf_2
Xhold553 _3853_/Q vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _3908_/Q vssd1 vssd1 vccd1 vccd1 _1902_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _3726_/Q vssd1 vssd1 vccd1 vccd1 _2702_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _3851_/Q vssd1 vssd1 vccd1 vccd1 _3177_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _4027_/Q vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold564 _3670_/X vssd1 vssd1 vccd1 vccd1 _4101_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _3506_/X _3507_/X _3508_/Y vssd1 vssd1 vccd1 vccd1 _3509_/X sky130_fd_sc_hd__a21o_1
Xhold586 _2838_/X vssd1 vssd1 vccd1 vccd1 _3780_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3213__A1 _3460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput40 _3808_/Q vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
Xoutput51 _3633_/A0 vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_12
XFILLER_0_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ _3860_/CLK _3860_/D vssd1 vssd1 vccd1 vccd1 _3860_/Q sky130_fd_sc_hd__dfxtp_1
X_3791_ _3791_/CLK _3791_/D vssd1 vssd1 vccd1 vccd1 _3791_/Q sky130_fd_sc_hd__dfxtp_1
X_2811_ _2869_/A _2811_/B _2813_/C vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__and3_1
XANTENNA__3204__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2742_ _3340_/A _2872_/A vssd1 vssd1 vccd1 vccd1 _2742_/X sky130_fd_sc_hd__and2_2
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2673_ _2813_/A _2673_/B _2676_/C vssd1 vssd1 vccd1 vccd1 _2673_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3225_ _3688_/Q _2681_/Y _3224_/X _3284_/A vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__o211a_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ hold292/X _3165_/B _3155_/X _3131_/A vssd1 vssd1 vccd1 vccd1 _3156_/X sky130_fd_sc_hd__o211a_1
X_3087_ _3171_/A _3133_/A vssd1 vssd1 vccd1 vccd1 _3087_/Y sky130_fd_sc_hd__nor2_1
X_2107_ _3905_/Q _3787_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2107_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2038_ _2034_/X _2037_/X _2119_/S vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _4112_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2113__S _2153_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 _3591_/X vssd1 vssd1 vccd1 vccd1 _4045_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _3211_/X vssd1 vssd1 vccd1 vccd1 _3867_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2182__B2 _2616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2182__A1 _1945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 _3742_/Q vssd1 vssd1 vccd1 vccd1 _2748_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _3761_/Q vssd1 vssd1 vccd1 vccd1 _2791_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _3357_/X vssd1 vssd1 vccd1 vccd1 _3936_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold479_A _3579_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2349__A _3518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2945__B1 _2953_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2023__S _2161_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3803_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3010_ _3060_/B _3008_/X _3009_/Y vssd1 vssd1 vccd1 vccd1 _3010_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3912_ _4101_/CLK _3912_/D vssd1 vssd1 vccd1 vccd1 _3912_/Q sky130_fd_sc_hd__dfxtp_1
X_3843_ _3846_/CLK _3843_/D vssd1 vssd1 vccd1 vccd1 _3843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3774_ _3791_/CLK _3774_/D vssd1 vssd1 vccd1 vccd1 _3774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2725_ _2887_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _3736_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2656_ _2652_/Y _2655_/X _2654_/X vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__a21o_1
X_2587_ _1880_/Y _2586_/X _2587_/S vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__mux2_1
Xfanout104 _2698_/A vssd1 vssd1 vccd1 vccd1 _2887_/A sky130_fd_sc_hd__clkbuf_4
X_3208_ _1889_/Y _3201_/A _2410_/B _2407_/A vssd1 vssd1 vccd1 vccd1 _3208_/X sky130_fd_sc_hd__a31o_1
X_3139_ hold326/X _3138_/A _3138_/Y _3320_/A vssd1 vssd1 vccd1 vccd1 _3139_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 _2601_/X vssd1 vssd1 vccd1 vccd1 _3701_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _3964_/Q vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2079__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3655__A1 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3402__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2018__S _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2510_ _2573_/S _3529_/A _2508_/Y _2509_/X vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__o22a_1
X_3490_ _1840_/A _3024_/A _3496_/S vssd1 vssd1 vccd1 vccd1 _3491_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2441_ _2585_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2441_/Y sky130_fd_sc_hd__nand2b_1
X_2372_ _2215_/C _2373_/B _2230_/B vssd1 vssd1 vccd1 vccd1 _2372_/Y sky130_fd_sc_hd__a21oi_1
X_4111_ _4111_/CLK _4111_/D vssd1 vssd1 vccd1 vccd1 _4111_/Q sky130_fd_sc_hd__dfxtp_1
X_4042_ _4042_/CLK _4042_/D vssd1 vssd1 vccd1 vccd1 _4042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3826_ _4077_/CLK _3826_/D vssd1 vssd1 vccd1 vccd1 _3826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ _3791_/CLK _3757_/D vssd1 vssd1 vccd1 vccd1 _3757_/Q sky130_fd_sc_hd__dfxtp_1
X_2708_ _3808_/Q _3247_/A vssd1 vssd1 vccd1 vccd1 _2708_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3688_ _4014_/CLK _3688_/D vssd1 vssd1 vccd1 vccd1 _3688_/Q sky130_fd_sc_hd__dfxtp_2
X_2639_ _3589_/A _2642_/B _2638_/Y _2734_/S _2164_/S vssd1 vssd1 vccd1 vccd1 _2639_/Y
+ sky130_fd_sc_hd__o32ai_1
XFILLER_0_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3458__A _3458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold609_A _3692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2679__A2 _2678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2990_ _3118_/B _3120_/A _2990_/C _2990_/D vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1941_ _2616_/B _1941_/B vssd1 vssd1 vccd1 vccd1 _2296_/C sky130_fd_sc_hd__nand2_1
X_1872_ _3829_/Q vssd1 vssd1 vccd1 vccd1 _3285_/B sky130_fd_sc_hd__inv_2
X_3611_ _3682_/A0 hold225/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3542_ _3529_/A _3525_/B _3541_/X vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3473_ hold581/X _3496_/S _3472_/Y _3587_/A vssd1 vssd1 vccd1 vccd1 _3473_/X sky130_fd_sc_hd__o211a_1
X_2424_ _2424_/A _2424_/B _2424_/C vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__and3_1
X_2355_ _1941_/B _2258_/Y _2354_/X vssd1 vssd1 vccd1 vccd1 _2355_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2286_ _2219_/B _4087_/Q vssd1 vssd1 vccd1 vccd1 _2288_/B sky130_fd_sc_hd__and2b_1
XANTENNA__3550__B _3551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _4031_/CLK _4025_/D vssd1 vssd1 vccd1 vccd1 _4025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3809_ _4111_/CLK _3809_/D vssd1 vssd1 vccd1 vccd1 _3809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2530__A1 _3637_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold559_A _3695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3188__A _3320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2444__S1 _2582_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _2138_/X _2139_/X _2158_/S vssd1 vssd1 vccd1 vccd1 _2140_/X sky130_fd_sc_hd__mux2_1
X_2071_ _3766_/Q _3750_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2071_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2973_ _3817_/Q _2971_/X hold606/X _3131_/A vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1924_ _2834_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _3323_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1855_ _3886_/Q vssd1 vssd1 vccd1 vccd1 _1855_/Y sky130_fd_sc_hd__inv_2
Xhold702 _3069_/X vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 _4083_/Q vssd1 vssd1 vccd1 vccd1 _3644_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold735 _3708_/Q vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _3130_/X vssd1 vssd1 vccd1 vccd1 _3131_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _4043_/Q vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ _3529_/A _3525_/B vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3456_ hold358/X _3676_/A0 _3470_/B vssd1 vssd1 vccd1 vccd1 _3456_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2407_ _2407_/A _2407_/B _2407_/C _2407_/D vssd1 vssd1 vccd1 vccd1 _2409_/A sky130_fd_sc_hd__or4_1
X_3387_ _3873_/Q _3874_/Q vssd1 vssd1 vccd1 vccd1 _3675_/A sky130_fd_sc_hd__nand2b_2
X_2338_ _2345_/S _2338_/B vssd1 vssd1 vccd1 vccd1 _2338_/X sky130_fd_sc_hd__or2_1
X_2269_ _2269_/A _2376_/B vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__or2_1
X_4008_ _4016_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2751__A1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2267__B1 _3554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_4 hold96/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3310_ hold657/X _3314_/S _3309_/X _3114_/A vssd1 vssd1 vccd1 vccd1 _3310_/X sky130_fd_sc_hd__o211a_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3587_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3886_/D sky130_fd_sc_hd__nand2_1
X_3172_ hold3/X _3189_/S _3320_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__a21o_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _3714_/Q _3726_/Q _2161_/S vssd1 vssd1 vccd1 vccd1 _2124_/B sky130_fd_sc_hd__mux2_1
X_2054_ _3775_/Q _3791_/Q _2159_/S vssd1 vssd1 vccd1 vccd1 _2054_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2725__A _2887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2956_ _3676_/A0 _2940_/X _2955_/Y vssd1 vssd1 vccd1 vccd1 _2956_/Y sky130_fd_sc_hd__a21oi_1
X_1907_ _3911_/Q _1996_/S vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__or2_1
X_2887_ _2887_/A _2887_/B _2887_/C vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__and3_1
X_1838_ _3658_/A vssd1 vssd1 vccd1 vccd1 _2009_/B sky130_fd_sc_hd__inv_2
Xhold510 _2753_/X vssd1 vssd1 vccd1 vccd1 _3744_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold554 _3181_/X vssd1 vssd1 vccd1 vccd1 _3182_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _3764_/Q vssd1 vssd1 vccd1 vccd1 _2799_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _3281_/X vssd1 vssd1 vccd1 vccd1 _3282_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _3685_/X vssd1 vssd1 vccd1 vccd1 _3872_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _3178_/X vssd1 vssd1 vccd1 vccd1 _3851_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _3889_/Q vssd1 vssd1 vccd1 vccd1 _1852_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _4099_/Q vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3506_/X _3507_/X _3554_/A vssd1 vssd1 vccd1 vccd1 _3508_/Y sky130_fd_sc_hd__o21ai_1
Xhold598 _3815_/Q vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_3439_ _3634_/A0 hold45/X _3444_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
XANTENNA__3291__A _3658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput52 _3634_/A0 vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
Xoutput30 _3639_/A0 vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
Xoutput41 _3835_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
XANTENNA__2488__B1 _3544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3405__S _3406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3790_ _3791_/CLK _3790_/D vssd1 vssd1 vccd1 vccd1 _3790_/Q sky130_fd_sc_hd__dfxtp_1
X_2810_ _2671_/X _2797_/X _2809_/X vssd1 vssd1 vccd1 vccd1 _3769_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2741_ _2740_/X _2655_/X _2741_/S vssd1 vssd1 vccd1 vccd1 _3739_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2672_ _2652_/Y _2671_/X _2669_/X vssd1 vssd1 vccd1 vccd1 _3714_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_78_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2715__B2 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3224_ _3224_/A _3224_/B vssd1 vssd1 vccd1 vccd1 _3224_/X sky130_fd_sc_hd__or2_1
.ends

